`timescale 1ns/1ps

module synapse_block_n #(
    parameter NUM_NEURONS  = 15,
    parameter PHASE_BITS   = 4,
    parameter WEIGHT_WIDTH = 5,
    parameter WEIGHT_FILE  = "weights2.hex"
)(
    input  wire [0:NUM_NEURONS-1] nout,
    output wire [0:NUM_NEURONS-1] nin
);

reg signed [4:0] w [0:14][0:14];

initial begin
        w[0][0] = 5'h00;
        w[0][1] = 5'h0C;
        w[0][2] = 5'h05;
        w[0][3] = 5'h04;
        w[0][4] = 5'h1C;
        w[0][5] = 5'h05;
        w[0][6] = 5'h0E;
        w[0][7] = 5'h05;
        w[0][8] = 5'h05;
        w[0][9] = 5'h0D;
        w[0][10] = 5'h1C;
        w[0][11] = 5'h1C;
        w[0][12] = 5'h0D;
        w[0][13] = 5'h0D;
        w[0][14] = 5'h02;
        w[1][0] = 5'h0C;
        w[1][1] = 5'h00;
        w[1][2] = 5'h04;
        w[1][3] = 5'h04;
        w[1][4] = 5'h1D;
        w[1][5] = 5'h03;
        w[1][6] = 5'h0C;
        w[1][7] = 5'h04;
        w[1][8] = 5'h04;
        w[1][9] = 5'h0D;
        w[1][10] = 5'h1D;
        w[1][11] = 5'h1C;
        w[1][12] = 5'h0C;
        w[1][13] = 5'h0C;
        w[1][14] = 5'h01;
        w[2][0] = 5'h05;
        w[2][1] = 5'h04;
        w[2][2] = 5'h00;
        w[2][3] = 5'h1C;
        w[2][4] = 5'h13;
        w[2][5] = 5'h0D;
        w[2][6] = 5'h05;
        w[2][7] = 5'h1B;
        w[2][8] = 5'h0C;
        w[2][9] = 5'h04;
        w[2][10] = 5'h13;
        w[2][11] = 5'h03;
        w[2][12] = 5'h04;
        w[2][13] = 5'h04;
        w[2][14] = 5'h0B;
        w[3][0] = 5'h04;
        w[3][1] = 5'h04;
        w[3][2] = 5'h1C;
        w[3][3] = 5'h00;
        w[3][4] = 5'h05;
        w[3][5] = 5'h1B;
        w[3][6] = 5'h05;
        w[3][7] = 5'h1C;
        w[3][8] = 5'h1C;
        w[3][9] = 5'h04;
        w[3][10] = 5'h05;
        w[3][11] = 5'h05;
        w[3][12] = 5'h03;
        w[3][13] = 5'h05;
        w[3][14] = 5'h1B;
        w[4][0] = 5'h1C;
        w[4][1] = 5'h1D;
        w[4][2] = 5'h13;
        w[4][3] = 5'h05;
        w[4][4] = 5'h00;
        w[4][5] = 5'h12;
        w[4][6] = 5'h1C;
        w[4][7] = 5'h05;
        w[4][8] = 5'h13;
        w[4][9] = 5'h1C;
        w[4][10] = 5'h0F;
        w[4][11] = 5'h1C;
        w[4][12] = 5'h1C;
        w[4][13] = 5'h1C;
        w[4][14] = 5'h13;
        w[5][0] = 5'h05;
        w[5][1] = 5'h03;
        w[5][2] = 5'h0D;
        w[5][3] = 5'h1B;
        w[5][4] = 5'h12;
        w[5][5] = 5'h00;
        w[5][6] = 5'h05;
        w[5][7] = 5'h1B;
        w[5][8] = 5'h0C;
        w[5][9] = 5'h04;
        w[5][10] = 5'h12;
        w[5][11] = 5'h03;
        w[5][12] = 5'h04;
        w[5][13] = 5'h04;
        w[5][14] = 5'h0C;
        w[6][0] = 5'h0E;
        w[6][1] = 5'h0C;
        w[6][2] = 5'h05;
        w[6][3] = 5'h05;
        w[6][4] = 5'h1C;
        w[6][5] = 5'h05;
        w[6][6] = 5'h00;
        w[6][7] = 5'h04;
        w[6][8] = 5'h05;
        w[6][9] = 5'h0D;
        w[6][10] = 5'h1C;
        w[6][11] = 5'h1D;
        w[6][12] = 5'h0D;
        w[6][13] = 5'h0E;
        w[6][14] = 5'h02;
        w[7][0] = 5'h05;
        w[7][1] = 5'h04;
        w[7][2] = 5'h1B;
        w[7][3] = 5'h1C;
        w[7][4] = 5'h05;
        w[7][5] = 5'h1B;
        w[7][6] = 5'h04;
        w[7][7] = 5'h00;
        w[7][8] = 5'h1D;
        w[7][9] = 5'h04;
        w[7][10] = 5'h05;
        w[7][11] = 5'h13;
        w[7][12] = 5'h05;
        w[7][13] = 5'h03;
        w[7][14] = 5'h1B;
        w[8][0] = 5'h05;
        w[8][1] = 5'h04;
        w[8][2] = 5'h0C;
        w[8][3] = 5'h1C;
        w[8][4] = 5'h13;
        w[8][5] = 5'h0C;
        w[8][6] = 5'h05;
        w[8][7] = 5'h1D;
        w[8][8] = 5'h00;
        w[8][9] = 5'h05;
        w[8][10] = 5'h13;
        w[8][11] = 5'h02;
        w[8][12] = 5'h05;
        w[8][13] = 5'h05;
        w[8][14] = 5'h0B;
        w[9][0] = 5'h0D;
        w[9][1] = 5'h0D;
        w[9][2] = 5'h04;
        w[9][3] = 5'h04;
        w[9][4] = 5'h1C;
        w[9][5] = 5'h04;
        w[9][6] = 5'h0D;
        w[9][7] = 5'h04;
        w[9][8] = 5'h05;
        w[9][9] = 5'h00;
        w[9][10] = 5'h1C;
        w[9][11] = 5'h1C;
        w[9][12] = 5'h0D;
        w[9][13] = 5'h0D;
        w[9][14] = 5'h02;
        w[10][0] = 5'h1C;
        w[10][1] = 5'h1D;
        w[10][2] = 5'h13;
        w[10][3] = 5'h05;
        w[10][4] = 5'h0F;
        w[10][5] = 5'h12;
        w[10][6] = 5'h1C;
        w[10][7] = 5'h05;
        w[10][8] = 5'h13;
        w[10][9] = 5'h1C;
        w[10][10] = 5'h00;
        w[10][11] = 5'h1C;
        w[10][12] = 5'h1C;
        w[10][13] = 5'h1C;
        w[10][14] = 5'h13;
        w[11][0] = 5'h1C;
        w[11][1] = 5'h1C;
        w[11][2] = 5'h03;
        w[11][3] = 5'h05;
        w[11][4] = 5'h1C;
        w[11][5] = 5'h03;
        w[11][6] = 5'h1D;
        w[11][7] = 5'h13;
        w[11][8] = 5'h02;
        w[11][9] = 5'h1C;
        w[11][10] = 5'h1C;
        w[11][11] = 5'h00;
        w[11][12] = 5'h1B;
        w[11][13] = 5'h1D;
        w[11][14] = 5'h04;
        w[12][0] = 5'h0D;
        w[12][1] = 5'h0C;
        w[12][2] = 5'h04;
        w[12][3] = 5'h03;
        w[12][4] = 5'h1C;
        w[12][5] = 5'h04;
        w[12][6] = 5'h0D;
        w[12][7] = 5'h05;
        w[12][8] = 5'h05;
        w[12][9] = 5'h0D;
        w[12][10] = 5'h1C;
        w[12][11] = 5'h1B;
        w[12][12] = 5'h00;
        w[12][13] = 5'h0D;
        w[12][14] = 5'h02;
        w[13][0] = 5'h0D;
        w[13][1] = 5'h0C;
        w[13][2] = 5'h04;
        w[13][3] = 5'h05;
        w[13][4] = 5'h1C;
        w[13][5] = 5'h04;
        w[13][6] = 5'h0E;
        w[13][7] = 5'h03;
        w[13][8] = 5'h05;
        w[13][9] = 5'h0D;
        w[13][10] = 5'h1C;
        w[13][11] = 5'h1D;
        w[13][12] = 5'h0D;
        w[13][13] = 5'h00;
        w[13][14] = 5'h03;
        w[14][0] = 5'h02;
        w[14][1] = 5'h01;
        w[14][2] = 5'h0B;
        w[14][3] = 5'h1B;
        w[14][4] = 5'h13;
        w[14][5] = 5'h0C;
        w[14][6] = 5'h02;
        w[14][7] = 5'h1B;
        w[14][8] = 5'h0B;
        w[14][9] = 5'h02;
        w[14][10] = 5'h13;
        w[14][11] = 5'h04;
        w[14][12] = 5'h02;
        w[14][13] = 5'h03;
        w[14][14] = 5'h00;
    end  

    // Generate block for parallel computation of each output n_in[i]
    genvar i, j;
    generate
        for (i = 0; i < 15; i = i + 1) begin : synapse_i
            // Array to hold individual terms: w[i][j] * n_out[j]
            wire signed [10:0] term [0:14];
            
            // Compute each term based on n_out[j]
            for (j = 0; j < 15; j = j + 1) begin : term_j
                assign term[j] = nout[j] ? w[i][j] : -w[i][j];
            end
            
            // Sum all terms combinatorially
            wire signed [10:0] sum = term[0] + term[1] + term[2] + term[3] + term[4] +
                                    term[5] + term[6] + term[7] + term[8] + term[9] +
                                    term[10] + term[11] + term[12] + term[13] + term[14];
            
            // Assign n_in[i] based on the sign of the sum
            
            assign nin[i] = (sum > 0) ? 1'b1 : 1'b0;
        end
    endgenerate

endmodule
