`timescale 1ns/1ps

module synapse_block_n #(
    parameter n  = 210
//    parameter PHASE_BITS   = 4,
//    parameter WEIGHT_WIDTH = 5,
//    parameter WEIGHT_FILE  = "weights2.hex"
)(
    input  wire [0:n-1] nout,
    output wire [0:n-1] nin
);

reg signed [4:0] w [0:n-1][0:n-1];
initial begin
w[0][0] = 5'b00000; w[0][1] = 5'b01111; w[0][2] = 5'b01111; w[0][3] = 5'b01111; w[0][4] = 5'b01111; w[0][5] = 5'b01111; w[0][6] = 5'b01111; w[0][7] = 5'b01111; w[0][8] = 5'b01111; w[0][9] = 5'b01111; w[0][10] = 5'b01111; w[0][11] = 5'b01111; w[0][12] = 5'b01111; w[0][13] = 5'b01111; w[0][14] = 5'b01111; w[0][15] = 5'b01111; w[0][16] = 5'b01111; w[0][17] = 5'b01111; w[0][18] = 5'b01111; w[0][19] = 5'b01111; w[0][20] = 5'b01111; w[0][21] = 5'b01111; w[0][22] = 5'b01111; w[0][23] = 5'b01111; w[0][24] = 5'b01111; w[0][25] = 5'b01111; w[0][26] = 5'b01111; w[0][27] = 5'b01111; w[0][28] = 5'b01111; w[0][29] = 5'b01111; w[0][30] = 5'b01111; w[0][31] = 5'b00000; w[0][32] = 5'b10000; w[0][33] = 5'b10000; w[0][34] = 5'b10000; w[0][35] = 5'b10000; w[0][36] = 5'b10000; w[0][37] = 5'b10000; w[0][38] = 5'b00000; w[0][39] = 5'b01111; w[0][40] = 5'b01111; w[0][41] = 5'b01111; w[0][42] = 5'b01111; w[0][43] = 5'b01111; w[0][44] = 5'b01111; w[0][45] = 5'b10000; w[0][46] = 5'b10000; w[0][47] = 5'b10000; w[0][48] = 5'b10000; w[0][49] = 5'b10000; w[0][50] = 5'b10000; w[0][51] = 5'b10000; w[0][52] = 5'b10000; w[0][53] = 5'b01111; w[0][54] = 5'b01111; w[0][55] = 5'b01111; w[0][56] = 5'b01111; w[0][57] = 5'b01111; w[0][58] = 5'b01111; w[0][59] = 5'b00000; w[0][60] = 5'b00000; w[0][61] = 5'b01111; w[0][62] = 5'b10000; w[0][63] = 5'b00000; w[0][64] = 5'b01111; w[0][65] = 5'b00000; w[0][66] = 5'b00000; w[0][67] = 5'b01111; w[0][68] = 5'b01111; w[0][69] = 5'b01111; w[0][70] = 5'b01111; w[0][71] = 5'b01111; w[0][72] = 5'b01111; w[0][73] = 5'b00000; w[0][74] = 5'b01111; w[0][75] = 5'b01111; w[0][76] = 5'b10000; w[0][77] = 5'b00000; w[0][78] = 5'b01111; w[0][79] = 5'b01111; w[0][80] = 5'b00000; w[0][81] = 5'b01111; w[0][82] = 5'b01111; w[0][83] = 5'b01111; w[0][84] = 5'b01111; w[0][85] = 5'b01111; w[0][86] = 5'b01111; w[0][87] = 5'b00000; w[0][88] = 5'b01111; w[0][89] = 5'b01111; w[0][90] = 5'b10000; w[0][91] = 5'b10000; w[0][92] = 5'b01111; w[0][93] = 5'b01111; w[0][94] = 5'b01111; w[0][95] = 5'b01111; w[0][96] = 5'b01111; w[0][97] = 5'b01111; w[0][98] = 5'b01111; w[0][99] = 5'b01111; w[0][100] = 5'b01111; w[0][101] = 5'b00000; w[0][102] = 5'b01111; w[0][103] = 5'b01111; w[0][104] = 5'b10000; w[0][105] = 5'b10000; w[0][106] = 5'b01111; w[0][107] = 5'b00000; w[0][108] = 5'b00000; w[0][109] = 5'b01111; w[0][110] = 5'b01111; w[0][111] = 5'b01111; w[0][112] = 5'b01111; w[0][113] = 5'b01111; w[0][114] = 5'b01111; w[0][115] = 5'b00000; w[0][116] = 5'b01111; w[0][117] = 5'b01111; w[0][118] = 5'b10000; w[0][119] = 5'b10000; w[0][120] = 5'b00000; w[0][121] = 5'b00000; w[0][122] = 5'b00000; w[0][123] = 5'b01111; w[0][124] = 5'b01111; w[0][125] = 5'b01111; w[0][126] = 5'b01111; w[0][127] = 5'b01111; w[0][128] = 5'b01111; w[0][129] = 5'b00000; w[0][130] = 5'b01111; w[0][131] = 5'b01111; w[0][132] = 5'b00000; w[0][133] = 5'b10000; w[0][134] = 5'b01111; w[0][135] = 5'b01111; w[0][136] = 5'b00000; w[0][137] = 5'b01111; w[0][138] = 5'b01111; w[0][139] = 5'b01111; w[0][140] = 5'b01111; w[0][141] = 5'b01111; w[0][142] = 5'b01111; w[0][143] = 5'b00000; w[0][144] = 5'b00000; w[0][145] = 5'b01111; w[0][146] = 5'b00000; w[0][147] = 5'b10000; w[0][148] = 5'b01111; w[0][149] = 5'b00000; w[0][150] = 5'b00000; w[0][151] = 5'b01111; w[0][152] = 5'b01111; w[0][153] = 5'b01111; w[0][154] = 5'b01111; w[0][155] = 5'b01111; w[0][156] = 5'b01111; w[0][157] = 5'b00000; w[0][158] = 5'b00000; w[0][159] = 5'b00000; w[0][160] = 5'b10000; w[0][161] = 5'b10000; w[0][162] = 5'b10000; w[0][163] = 5'b00000; w[0][164] = 5'b00000; w[0][165] = 5'b01111; w[0][166] = 5'b01111; w[0][167] = 5'b01111; w[0][168] = 5'b01111; w[0][169] = 5'b01111; w[0][170] = 5'b01111; w[0][171] = 5'b01111; w[0][172] = 5'b00000; w[0][173] = 5'b00000; w[0][174] = 5'b10000; w[0][175] = 5'b10000; w[0][176] = 5'b10000; w[0][177] = 5'b00000; w[0][178] = 5'b01111; w[0][179] = 5'b01111; w[0][180] = 5'b01111; w[0][181] = 5'b01111; w[0][182] = 5'b01111; w[0][183] = 5'b01111; w[0][184] = 5'b01111; w[0][185] = 5'b01111; w[0][186] = 5'b01111; w[0][187] = 5'b01111; w[0][188] = 5'b01111; w[0][189] = 5'b01111; w[0][190] = 5'b01111; w[0][191] = 5'b01111; w[0][192] = 5'b01111; w[0][193] = 5'b01111; w[0][194] = 5'b01111; w[0][195] = 5'b01111; w[0][196] = 5'b01111; w[0][197] = 5'b01111; w[0][198] = 5'b01111; w[0][199] = 5'b01111; w[0][200] = 5'b01111; w[0][201] = 5'b01111; w[0][202] = 5'b01111; w[0][203] = 5'b01111; w[0][204] = 5'b01111; w[0][205] = 5'b01111; w[0][206] = 5'b01111; w[0][207] = 5'b01111; w[0][208] = 5'b01111; w[0][209] = 5'b01111; 
w[1][0] = 5'b01111; w[1][1] = 5'b00000; w[1][2] = 5'b01111; w[1][3] = 5'b01111; w[1][4] = 5'b01111; w[1][5] = 5'b01111; w[1][6] = 5'b01111; w[1][7] = 5'b01111; w[1][8] = 5'b01111; w[1][9] = 5'b01111; w[1][10] = 5'b01111; w[1][11] = 5'b01111; w[1][12] = 5'b01111; w[1][13] = 5'b01111; w[1][14] = 5'b01111; w[1][15] = 5'b01111; w[1][16] = 5'b01111; w[1][17] = 5'b01111; w[1][18] = 5'b01111; w[1][19] = 5'b01111; w[1][20] = 5'b01111; w[1][21] = 5'b01111; w[1][22] = 5'b01111; w[1][23] = 5'b01111; w[1][24] = 5'b01111; w[1][25] = 5'b01111; w[1][26] = 5'b01111; w[1][27] = 5'b01111; w[1][28] = 5'b01111; w[1][29] = 5'b01111; w[1][30] = 5'b01111; w[1][31] = 5'b00000; w[1][32] = 5'b10000; w[1][33] = 5'b10000; w[1][34] = 5'b10000; w[1][35] = 5'b10000; w[1][36] = 5'b10000; w[1][37] = 5'b10000; w[1][38] = 5'b00000; w[1][39] = 5'b01111; w[1][40] = 5'b01111; w[1][41] = 5'b01111; w[1][42] = 5'b01111; w[1][43] = 5'b01111; w[1][44] = 5'b01111; w[1][45] = 5'b10000; w[1][46] = 5'b10000; w[1][47] = 5'b10000; w[1][48] = 5'b10000; w[1][49] = 5'b10000; w[1][50] = 5'b10000; w[1][51] = 5'b10000; w[1][52] = 5'b10000; w[1][53] = 5'b01111; w[1][54] = 5'b01111; w[1][55] = 5'b01111; w[1][56] = 5'b01111; w[1][57] = 5'b01111; w[1][58] = 5'b01111; w[1][59] = 5'b00000; w[1][60] = 5'b00000; w[1][61] = 5'b01111; w[1][62] = 5'b10000; w[1][63] = 5'b00000; w[1][64] = 5'b01111; w[1][65] = 5'b00000; w[1][66] = 5'b00000; w[1][67] = 5'b01111; w[1][68] = 5'b01111; w[1][69] = 5'b01111; w[1][70] = 5'b01111; w[1][71] = 5'b01111; w[1][72] = 5'b01111; w[1][73] = 5'b00000; w[1][74] = 5'b01111; w[1][75] = 5'b01111; w[1][76] = 5'b10000; w[1][77] = 5'b00000; w[1][78] = 5'b01111; w[1][79] = 5'b01111; w[1][80] = 5'b00000; w[1][81] = 5'b01111; w[1][82] = 5'b01111; w[1][83] = 5'b01111; w[1][84] = 5'b01111; w[1][85] = 5'b01111; w[1][86] = 5'b01111; w[1][87] = 5'b00000; w[1][88] = 5'b01111; w[1][89] = 5'b01111; w[1][90] = 5'b10000; w[1][91] = 5'b10000; w[1][92] = 5'b01111; w[1][93] = 5'b01111; w[1][94] = 5'b01111; w[1][95] = 5'b01111; w[1][96] = 5'b01111; w[1][97] = 5'b01111; w[1][98] = 5'b01111; w[1][99] = 5'b01111; w[1][100] = 5'b01111; w[1][101] = 5'b00000; w[1][102] = 5'b01111; w[1][103] = 5'b01111; w[1][104] = 5'b10000; w[1][105] = 5'b10000; w[1][106] = 5'b01111; w[1][107] = 5'b00000; w[1][108] = 5'b00000; w[1][109] = 5'b01111; w[1][110] = 5'b01111; w[1][111] = 5'b01111; w[1][112] = 5'b01111; w[1][113] = 5'b01111; w[1][114] = 5'b01111; w[1][115] = 5'b00000; w[1][116] = 5'b01111; w[1][117] = 5'b01111; w[1][118] = 5'b10000; w[1][119] = 5'b10000; w[1][120] = 5'b00000; w[1][121] = 5'b00000; w[1][122] = 5'b00000; w[1][123] = 5'b01111; w[1][124] = 5'b01111; w[1][125] = 5'b01111; w[1][126] = 5'b01111; w[1][127] = 5'b01111; w[1][128] = 5'b01111; w[1][129] = 5'b00000; w[1][130] = 5'b01111; w[1][131] = 5'b01111; w[1][132] = 5'b00000; w[1][133] = 5'b10000; w[1][134] = 5'b01111; w[1][135] = 5'b01111; w[1][136] = 5'b00000; w[1][137] = 5'b01111; w[1][138] = 5'b01111; w[1][139] = 5'b01111; w[1][140] = 5'b01111; w[1][141] = 5'b01111; w[1][142] = 5'b01111; w[1][143] = 5'b00000; w[1][144] = 5'b00000; w[1][145] = 5'b01111; w[1][146] = 5'b00000; w[1][147] = 5'b10000; w[1][148] = 5'b01111; w[1][149] = 5'b00000; w[1][150] = 5'b00000; w[1][151] = 5'b01111; w[1][152] = 5'b01111; w[1][153] = 5'b01111; w[1][154] = 5'b01111; w[1][155] = 5'b01111; w[1][156] = 5'b01111; w[1][157] = 5'b00000; w[1][158] = 5'b00000; w[1][159] = 5'b00000; w[1][160] = 5'b10000; w[1][161] = 5'b10000; w[1][162] = 5'b10000; w[1][163] = 5'b00000; w[1][164] = 5'b00000; w[1][165] = 5'b01111; w[1][166] = 5'b01111; w[1][167] = 5'b01111; w[1][168] = 5'b01111; w[1][169] = 5'b01111; w[1][170] = 5'b01111; w[1][171] = 5'b01111; w[1][172] = 5'b00000; w[1][173] = 5'b00000; w[1][174] = 5'b10000; w[1][175] = 5'b10000; w[1][176] = 5'b10000; w[1][177] = 5'b00000; w[1][178] = 5'b01111; w[1][179] = 5'b01111; w[1][180] = 5'b01111; w[1][181] = 5'b01111; w[1][182] = 5'b01111; w[1][183] = 5'b01111; w[1][184] = 5'b01111; w[1][185] = 5'b01111; w[1][186] = 5'b01111; w[1][187] = 5'b01111; w[1][188] = 5'b01111; w[1][189] = 5'b01111; w[1][190] = 5'b01111; w[1][191] = 5'b01111; w[1][192] = 5'b01111; w[1][193] = 5'b01111; w[1][194] = 5'b01111; w[1][195] = 5'b01111; w[1][196] = 5'b01111; w[1][197] = 5'b01111; w[1][198] = 5'b01111; w[1][199] = 5'b01111; w[1][200] = 5'b01111; w[1][201] = 5'b01111; w[1][202] = 5'b01111; w[1][203] = 5'b01111; w[1][204] = 5'b01111; w[1][205] = 5'b01111; w[1][206] = 5'b01111; w[1][207] = 5'b01111; w[1][208] = 5'b01111; w[1][209] = 5'b01111; 
w[2][0] = 5'b01111; w[2][1] = 5'b01111; w[2][2] = 5'b00000; w[2][3] = 5'b01111; w[2][4] = 5'b01111; w[2][5] = 5'b01111; w[2][6] = 5'b01111; w[2][7] = 5'b01111; w[2][8] = 5'b01111; w[2][9] = 5'b01111; w[2][10] = 5'b01111; w[2][11] = 5'b01111; w[2][12] = 5'b01111; w[2][13] = 5'b01111; w[2][14] = 5'b01111; w[2][15] = 5'b01111; w[2][16] = 5'b01111; w[2][17] = 5'b01111; w[2][18] = 5'b01111; w[2][19] = 5'b01111; w[2][20] = 5'b01111; w[2][21] = 5'b01111; w[2][22] = 5'b01111; w[2][23] = 5'b01111; w[2][24] = 5'b01111; w[2][25] = 5'b01111; w[2][26] = 5'b01111; w[2][27] = 5'b01111; w[2][28] = 5'b01111; w[2][29] = 5'b01111; w[2][30] = 5'b01111; w[2][31] = 5'b00000; w[2][32] = 5'b10000; w[2][33] = 5'b10000; w[2][34] = 5'b10000; w[2][35] = 5'b10000; w[2][36] = 5'b10000; w[2][37] = 5'b10000; w[2][38] = 5'b00000; w[2][39] = 5'b01111; w[2][40] = 5'b01111; w[2][41] = 5'b01111; w[2][42] = 5'b01111; w[2][43] = 5'b01111; w[2][44] = 5'b01111; w[2][45] = 5'b10000; w[2][46] = 5'b10000; w[2][47] = 5'b10000; w[2][48] = 5'b10000; w[2][49] = 5'b10000; w[2][50] = 5'b10000; w[2][51] = 5'b10000; w[2][52] = 5'b10000; w[2][53] = 5'b01111; w[2][54] = 5'b01111; w[2][55] = 5'b01111; w[2][56] = 5'b01111; w[2][57] = 5'b01111; w[2][58] = 5'b01111; w[2][59] = 5'b00000; w[2][60] = 5'b00000; w[2][61] = 5'b01111; w[2][62] = 5'b10000; w[2][63] = 5'b00000; w[2][64] = 5'b01111; w[2][65] = 5'b00000; w[2][66] = 5'b00000; w[2][67] = 5'b01111; w[2][68] = 5'b01111; w[2][69] = 5'b01111; w[2][70] = 5'b01111; w[2][71] = 5'b01111; w[2][72] = 5'b01111; w[2][73] = 5'b00000; w[2][74] = 5'b01111; w[2][75] = 5'b01111; w[2][76] = 5'b10000; w[2][77] = 5'b00000; w[2][78] = 5'b01111; w[2][79] = 5'b01111; w[2][80] = 5'b00000; w[2][81] = 5'b01111; w[2][82] = 5'b01111; w[2][83] = 5'b01111; w[2][84] = 5'b01111; w[2][85] = 5'b01111; w[2][86] = 5'b01111; w[2][87] = 5'b00000; w[2][88] = 5'b01111; w[2][89] = 5'b01111; w[2][90] = 5'b10000; w[2][91] = 5'b10000; w[2][92] = 5'b01111; w[2][93] = 5'b01111; w[2][94] = 5'b01111; w[2][95] = 5'b01111; w[2][96] = 5'b01111; w[2][97] = 5'b01111; w[2][98] = 5'b01111; w[2][99] = 5'b01111; w[2][100] = 5'b01111; w[2][101] = 5'b00000; w[2][102] = 5'b01111; w[2][103] = 5'b01111; w[2][104] = 5'b10000; w[2][105] = 5'b10000; w[2][106] = 5'b01111; w[2][107] = 5'b00000; w[2][108] = 5'b00000; w[2][109] = 5'b01111; w[2][110] = 5'b01111; w[2][111] = 5'b01111; w[2][112] = 5'b01111; w[2][113] = 5'b01111; w[2][114] = 5'b01111; w[2][115] = 5'b00000; w[2][116] = 5'b01111; w[2][117] = 5'b01111; w[2][118] = 5'b10000; w[2][119] = 5'b10000; w[2][120] = 5'b00000; w[2][121] = 5'b00000; w[2][122] = 5'b00000; w[2][123] = 5'b01111; w[2][124] = 5'b01111; w[2][125] = 5'b01111; w[2][126] = 5'b01111; w[2][127] = 5'b01111; w[2][128] = 5'b01111; w[2][129] = 5'b00000; w[2][130] = 5'b01111; w[2][131] = 5'b01111; w[2][132] = 5'b00000; w[2][133] = 5'b10000; w[2][134] = 5'b01111; w[2][135] = 5'b01111; w[2][136] = 5'b00000; w[2][137] = 5'b01111; w[2][138] = 5'b01111; w[2][139] = 5'b01111; w[2][140] = 5'b01111; w[2][141] = 5'b01111; w[2][142] = 5'b01111; w[2][143] = 5'b00000; w[2][144] = 5'b00000; w[2][145] = 5'b01111; w[2][146] = 5'b00000; w[2][147] = 5'b10000; w[2][148] = 5'b01111; w[2][149] = 5'b00000; w[2][150] = 5'b00000; w[2][151] = 5'b01111; w[2][152] = 5'b01111; w[2][153] = 5'b01111; w[2][154] = 5'b01111; w[2][155] = 5'b01111; w[2][156] = 5'b01111; w[2][157] = 5'b00000; w[2][158] = 5'b00000; w[2][159] = 5'b00000; w[2][160] = 5'b10000; w[2][161] = 5'b10000; w[2][162] = 5'b10000; w[2][163] = 5'b00000; w[2][164] = 5'b00000; w[2][165] = 5'b01111; w[2][166] = 5'b01111; w[2][167] = 5'b01111; w[2][168] = 5'b01111; w[2][169] = 5'b01111; w[2][170] = 5'b01111; w[2][171] = 5'b01111; w[2][172] = 5'b00000; w[2][173] = 5'b00000; w[2][174] = 5'b10000; w[2][175] = 5'b10000; w[2][176] = 5'b10000; w[2][177] = 5'b00000; w[2][178] = 5'b01111; w[2][179] = 5'b01111; w[2][180] = 5'b01111; w[2][181] = 5'b01111; w[2][182] = 5'b01111; w[2][183] = 5'b01111; w[2][184] = 5'b01111; w[2][185] = 5'b01111; w[2][186] = 5'b01111; w[2][187] = 5'b01111; w[2][188] = 5'b01111; w[2][189] = 5'b01111; w[2][190] = 5'b01111; w[2][191] = 5'b01111; w[2][192] = 5'b01111; w[2][193] = 5'b01111; w[2][194] = 5'b01111; w[2][195] = 5'b01111; w[2][196] = 5'b01111; w[2][197] = 5'b01111; w[2][198] = 5'b01111; w[2][199] = 5'b01111; w[2][200] = 5'b01111; w[2][201] = 5'b01111; w[2][202] = 5'b01111; w[2][203] = 5'b01111; w[2][204] = 5'b01111; w[2][205] = 5'b01111; w[2][206] = 5'b01111; w[2][207] = 5'b01111; w[2][208] = 5'b01111; w[2][209] = 5'b01111; 
w[3][0] = 5'b01111; w[3][1] = 5'b01111; w[3][2] = 5'b01111; w[3][3] = 5'b00000; w[3][4] = 5'b01111; w[3][5] = 5'b01111; w[3][6] = 5'b01111; w[3][7] = 5'b01111; w[3][8] = 5'b01111; w[3][9] = 5'b01111; w[3][10] = 5'b01111; w[3][11] = 5'b01111; w[3][12] = 5'b01111; w[3][13] = 5'b01111; w[3][14] = 5'b01111; w[3][15] = 5'b01111; w[3][16] = 5'b01111; w[3][17] = 5'b01111; w[3][18] = 5'b01111; w[3][19] = 5'b01111; w[3][20] = 5'b01111; w[3][21] = 5'b01111; w[3][22] = 5'b01111; w[3][23] = 5'b01111; w[3][24] = 5'b01111; w[3][25] = 5'b01111; w[3][26] = 5'b01111; w[3][27] = 5'b01111; w[3][28] = 5'b01111; w[3][29] = 5'b01111; w[3][30] = 5'b01111; w[3][31] = 5'b00000; w[3][32] = 5'b10000; w[3][33] = 5'b10000; w[3][34] = 5'b10000; w[3][35] = 5'b10000; w[3][36] = 5'b10000; w[3][37] = 5'b10000; w[3][38] = 5'b00000; w[3][39] = 5'b01111; w[3][40] = 5'b01111; w[3][41] = 5'b01111; w[3][42] = 5'b01111; w[3][43] = 5'b01111; w[3][44] = 5'b01111; w[3][45] = 5'b10000; w[3][46] = 5'b10000; w[3][47] = 5'b10000; w[3][48] = 5'b10000; w[3][49] = 5'b10000; w[3][50] = 5'b10000; w[3][51] = 5'b10000; w[3][52] = 5'b10000; w[3][53] = 5'b01111; w[3][54] = 5'b01111; w[3][55] = 5'b01111; w[3][56] = 5'b01111; w[3][57] = 5'b01111; w[3][58] = 5'b01111; w[3][59] = 5'b00000; w[3][60] = 5'b00000; w[3][61] = 5'b01111; w[3][62] = 5'b10000; w[3][63] = 5'b00000; w[3][64] = 5'b01111; w[3][65] = 5'b00000; w[3][66] = 5'b00000; w[3][67] = 5'b01111; w[3][68] = 5'b01111; w[3][69] = 5'b01111; w[3][70] = 5'b01111; w[3][71] = 5'b01111; w[3][72] = 5'b01111; w[3][73] = 5'b00000; w[3][74] = 5'b01111; w[3][75] = 5'b01111; w[3][76] = 5'b10000; w[3][77] = 5'b00000; w[3][78] = 5'b01111; w[3][79] = 5'b01111; w[3][80] = 5'b00000; w[3][81] = 5'b01111; w[3][82] = 5'b01111; w[3][83] = 5'b01111; w[3][84] = 5'b01111; w[3][85] = 5'b01111; w[3][86] = 5'b01111; w[3][87] = 5'b00000; w[3][88] = 5'b01111; w[3][89] = 5'b01111; w[3][90] = 5'b10000; w[3][91] = 5'b10000; w[3][92] = 5'b01111; w[3][93] = 5'b01111; w[3][94] = 5'b01111; w[3][95] = 5'b01111; w[3][96] = 5'b01111; w[3][97] = 5'b01111; w[3][98] = 5'b01111; w[3][99] = 5'b01111; w[3][100] = 5'b01111; w[3][101] = 5'b00000; w[3][102] = 5'b01111; w[3][103] = 5'b01111; w[3][104] = 5'b10000; w[3][105] = 5'b10000; w[3][106] = 5'b01111; w[3][107] = 5'b00000; w[3][108] = 5'b00000; w[3][109] = 5'b01111; w[3][110] = 5'b01111; w[3][111] = 5'b01111; w[3][112] = 5'b01111; w[3][113] = 5'b01111; w[3][114] = 5'b01111; w[3][115] = 5'b00000; w[3][116] = 5'b01111; w[3][117] = 5'b01111; w[3][118] = 5'b10000; w[3][119] = 5'b10000; w[3][120] = 5'b00000; w[3][121] = 5'b00000; w[3][122] = 5'b00000; w[3][123] = 5'b01111; w[3][124] = 5'b01111; w[3][125] = 5'b01111; w[3][126] = 5'b01111; w[3][127] = 5'b01111; w[3][128] = 5'b01111; w[3][129] = 5'b00000; w[3][130] = 5'b01111; w[3][131] = 5'b01111; w[3][132] = 5'b00000; w[3][133] = 5'b10000; w[3][134] = 5'b01111; w[3][135] = 5'b01111; w[3][136] = 5'b00000; w[3][137] = 5'b01111; w[3][138] = 5'b01111; w[3][139] = 5'b01111; w[3][140] = 5'b01111; w[3][141] = 5'b01111; w[3][142] = 5'b01111; w[3][143] = 5'b00000; w[3][144] = 5'b00000; w[3][145] = 5'b01111; w[3][146] = 5'b00000; w[3][147] = 5'b10000; w[3][148] = 5'b01111; w[3][149] = 5'b00000; w[3][150] = 5'b00000; w[3][151] = 5'b01111; w[3][152] = 5'b01111; w[3][153] = 5'b01111; w[3][154] = 5'b01111; w[3][155] = 5'b01111; w[3][156] = 5'b01111; w[3][157] = 5'b00000; w[3][158] = 5'b00000; w[3][159] = 5'b00000; w[3][160] = 5'b10000; w[3][161] = 5'b10000; w[3][162] = 5'b10000; w[3][163] = 5'b00000; w[3][164] = 5'b00000; w[3][165] = 5'b01111; w[3][166] = 5'b01111; w[3][167] = 5'b01111; w[3][168] = 5'b01111; w[3][169] = 5'b01111; w[3][170] = 5'b01111; w[3][171] = 5'b01111; w[3][172] = 5'b00000; w[3][173] = 5'b00000; w[3][174] = 5'b10000; w[3][175] = 5'b10000; w[3][176] = 5'b10000; w[3][177] = 5'b00000; w[3][178] = 5'b01111; w[3][179] = 5'b01111; w[3][180] = 5'b01111; w[3][181] = 5'b01111; w[3][182] = 5'b01111; w[3][183] = 5'b01111; w[3][184] = 5'b01111; w[3][185] = 5'b01111; w[3][186] = 5'b01111; w[3][187] = 5'b01111; w[3][188] = 5'b01111; w[3][189] = 5'b01111; w[3][190] = 5'b01111; w[3][191] = 5'b01111; w[3][192] = 5'b01111; w[3][193] = 5'b01111; w[3][194] = 5'b01111; w[3][195] = 5'b01111; w[3][196] = 5'b01111; w[3][197] = 5'b01111; w[3][198] = 5'b01111; w[3][199] = 5'b01111; w[3][200] = 5'b01111; w[3][201] = 5'b01111; w[3][202] = 5'b01111; w[3][203] = 5'b01111; w[3][204] = 5'b01111; w[3][205] = 5'b01111; w[3][206] = 5'b01111; w[3][207] = 5'b01111; w[3][208] = 5'b01111; w[3][209] = 5'b01111; 
w[4][0] = 5'b01111; w[4][1] = 5'b01111; w[4][2] = 5'b01111; w[4][3] = 5'b01111; w[4][4] = 5'b00000; w[4][5] = 5'b01111; w[4][6] = 5'b01111; w[4][7] = 5'b01111; w[4][8] = 5'b01111; w[4][9] = 5'b01111; w[4][10] = 5'b01111; w[4][11] = 5'b01111; w[4][12] = 5'b01111; w[4][13] = 5'b01111; w[4][14] = 5'b01111; w[4][15] = 5'b01111; w[4][16] = 5'b01111; w[4][17] = 5'b01111; w[4][18] = 5'b01111; w[4][19] = 5'b01111; w[4][20] = 5'b01111; w[4][21] = 5'b01111; w[4][22] = 5'b01111; w[4][23] = 5'b01111; w[4][24] = 5'b01111; w[4][25] = 5'b01111; w[4][26] = 5'b01111; w[4][27] = 5'b01111; w[4][28] = 5'b01111; w[4][29] = 5'b01111; w[4][30] = 5'b01111; w[4][31] = 5'b00000; w[4][32] = 5'b10000; w[4][33] = 5'b10000; w[4][34] = 5'b10000; w[4][35] = 5'b10000; w[4][36] = 5'b10000; w[4][37] = 5'b10000; w[4][38] = 5'b00000; w[4][39] = 5'b01111; w[4][40] = 5'b01111; w[4][41] = 5'b01111; w[4][42] = 5'b01111; w[4][43] = 5'b01111; w[4][44] = 5'b01111; w[4][45] = 5'b10000; w[4][46] = 5'b10000; w[4][47] = 5'b10000; w[4][48] = 5'b10000; w[4][49] = 5'b10000; w[4][50] = 5'b10000; w[4][51] = 5'b10000; w[4][52] = 5'b10000; w[4][53] = 5'b01111; w[4][54] = 5'b01111; w[4][55] = 5'b01111; w[4][56] = 5'b01111; w[4][57] = 5'b01111; w[4][58] = 5'b01111; w[4][59] = 5'b00000; w[4][60] = 5'b00000; w[4][61] = 5'b01111; w[4][62] = 5'b10000; w[4][63] = 5'b00000; w[4][64] = 5'b01111; w[4][65] = 5'b00000; w[4][66] = 5'b00000; w[4][67] = 5'b01111; w[4][68] = 5'b01111; w[4][69] = 5'b01111; w[4][70] = 5'b01111; w[4][71] = 5'b01111; w[4][72] = 5'b01111; w[4][73] = 5'b00000; w[4][74] = 5'b01111; w[4][75] = 5'b01111; w[4][76] = 5'b10000; w[4][77] = 5'b00000; w[4][78] = 5'b01111; w[4][79] = 5'b01111; w[4][80] = 5'b00000; w[4][81] = 5'b01111; w[4][82] = 5'b01111; w[4][83] = 5'b01111; w[4][84] = 5'b01111; w[4][85] = 5'b01111; w[4][86] = 5'b01111; w[4][87] = 5'b00000; w[4][88] = 5'b01111; w[4][89] = 5'b01111; w[4][90] = 5'b10000; w[4][91] = 5'b10000; w[4][92] = 5'b01111; w[4][93] = 5'b01111; w[4][94] = 5'b01111; w[4][95] = 5'b01111; w[4][96] = 5'b01111; w[4][97] = 5'b01111; w[4][98] = 5'b01111; w[4][99] = 5'b01111; w[4][100] = 5'b01111; w[4][101] = 5'b00000; w[4][102] = 5'b01111; w[4][103] = 5'b01111; w[4][104] = 5'b10000; w[4][105] = 5'b10000; w[4][106] = 5'b01111; w[4][107] = 5'b00000; w[4][108] = 5'b00000; w[4][109] = 5'b01111; w[4][110] = 5'b01111; w[4][111] = 5'b01111; w[4][112] = 5'b01111; w[4][113] = 5'b01111; w[4][114] = 5'b01111; w[4][115] = 5'b00000; w[4][116] = 5'b01111; w[4][117] = 5'b01111; w[4][118] = 5'b10000; w[4][119] = 5'b10000; w[4][120] = 5'b00000; w[4][121] = 5'b00000; w[4][122] = 5'b00000; w[4][123] = 5'b01111; w[4][124] = 5'b01111; w[4][125] = 5'b01111; w[4][126] = 5'b01111; w[4][127] = 5'b01111; w[4][128] = 5'b01111; w[4][129] = 5'b00000; w[4][130] = 5'b01111; w[4][131] = 5'b01111; w[4][132] = 5'b00000; w[4][133] = 5'b10000; w[4][134] = 5'b01111; w[4][135] = 5'b01111; w[4][136] = 5'b00000; w[4][137] = 5'b01111; w[4][138] = 5'b01111; w[4][139] = 5'b01111; w[4][140] = 5'b01111; w[4][141] = 5'b01111; w[4][142] = 5'b01111; w[4][143] = 5'b00000; w[4][144] = 5'b00000; w[4][145] = 5'b01111; w[4][146] = 5'b00000; w[4][147] = 5'b10000; w[4][148] = 5'b01111; w[4][149] = 5'b00000; w[4][150] = 5'b00000; w[4][151] = 5'b01111; w[4][152] = 5'b01111; w[4][153] = 5'b01111; w[4][154] = 5'b01111; w[4][155] = 5'b01111; w[4][156] = 5'b01111; w[4][157] = 5'b00000; w[4][158] = 5'b00000; w[4][159] = 5'b00000; w[4][160] = 5'b10000; w[4][161] = 5'b10000; w[4][162] = 5'b10000; w[4][163] = 5'b00000; w[4][164] = 5'b00000; w[4][165] = 5'b01111; w[4][166] = 5'b01111; w[4][167] = 5'b01111; w[4][168] = 5'b01111; w[4][169] = 5'b01111; w[4][170] = 5'b01111; w[4][171] = 5'b01111; w[4][172] = 5'b00000; w[4][173] = 5'b00000; w[4][174] = 5'b10000; w[4][175] = 5'b10000; w[4][176] = 5'b10000; w[4][177] = 5'b00000; w[4][178] = 5'b01111; w[4][179] = 5'b01111; w[4][180] = 5'b01111; w[4][181] = 5'b01111; w[4][182] = 5'b01111; w[4][183] = 5'b01111; w[4][184] = 5'b01111; w[4][185] = 5'b01111; w[4][186] = 5'b01111; w[4][187] = 5'b01111; w[4][188] = 5'b01111; w[4][189] = 5'b01111; w[4][190] = 5'b01111; w[4][191] = 5'b01111; w[4][192] = 5'b01111; w[4][193] = 5'b01111; w[4][194] = 5'b01111; w[4][195] = 5'b01111; w[4][196] = 5'b01111; w[4][197] = 5'b01111; w[4][198] = 5'b01111; w[4][199] = 5'b01111; w[4][200] = 5'b01111; w[4][201] = 5'b01111; w[4][202] = 5'b01111; w[4][203] = 5'b01111; w[4][204] = 5'b01111; w[4][205] = 5'b01111; w[4][206] = 5'b01111; w[4][207] = 5'b01111; w[4][208] = 5'b01111; w[4][209] = 5'b01111; 
w[5][0] = 5'b01111; w[5][1] = 5'b01111; w[5][2] = 5'b01111; w[5][3] = 5'b01111; w[5][4] = 5'b01111; w[5][5] = 5'b00000; w[5][6] = 5'b01111; w[5][7] = 5'b01111; w[5][8] = 5'b01111; w[5][9] = 5'b01111; w[5][10] = 5'b01111; w[5][11] = 5'b01111; w[5][12] = 5'b01111; w[5][13] = 5'b01111; w[5][14] = 5'b01111; w[5][15] = 5'b01111; w[5][16] = 5'b01111; w[5][17] = 5'b01111; w[5][18] = 5'b01111; w[5][19] = 5'b01111; w[5][20] = 5'b01111; w[5][21] = 5'b01111; w[5][22] = 5'b01111; w[5][23] = 5'b01111; w[5][24] = 5'b01111; w[5][25] = 5'b01111; w[5][26] = 5'b01111; w[5][27] = 5'b01111; w[5][28] = 5'b01111; w[5][29] = 5'b01111; w[5][30] = 5'b01111; w[5][31] = 5'b00000; w[5][32] = 5'b10000; w[5][33] = 5'b10000; w[5][34] = 5'b10000; w[5][35] = 5'b10000; w[5][36] = 5'b10000; w[5][37] = 5'b10000; w[5][38] = 5'b00000; w[5][39] = 5'b01111; w[5][40] = 5'b01111; w[5][41] = 5'b01111; w[5][42] = 5'b01111; w[5][43] = 5'b01111; w[5][44] = 5'b01111; w[5][45] = 5'b10000; w[5][46] = 5'b10000; w[5][47] = 5'b10000; w[5][48] = 5'b10000; w[5][49] = 5'b10000; w[5][50] = 5'b10000; w[5][51] = 5'b10000; w[5][52] = 5'b10000; w[5][53] = 5'b01111; w[5][54] = 5'b01111; w[5][55] = 5'b01111; w[5][56] = 5'b01111; w[5][57] = 5'b01111; w[5][58] = 5'b01111; w[5][59] = 5'b00000; w[5][60] = 5'b00000; w[5][61] = 5'b01111; w[5][62] = 5'b10000; w[5][63] = 5'b00000; w[5][64] = 5'b01111; w[5][65] = 5'b00000; w[5][66] = 5'b00000; w[5][67] = 5'b01111; w[5][68] = 5'b01111; w[5][69] = 5'b01111; w[5][70] = 5'b01111; w[5][71] = 5'b01111; w[5][72] = 5'b01111; w[5][73] = 5'b00000; w[5][74] = 5'b01111; w[5][75] = 5'b01111; w[5][76] = 5'b10000; w[5][77] = 5'b00000; w[5][78] = 5'b01111; w[5][79] = 5'b01111; w[5][80] = 5'b00000; w[5][81] = 5'b01111; w[5][82] = 5'b01111; w[5][83] = 5'b01111; w[5][84] = 5'b01111; w[5][85] = 5'b01111; w[5][86] = 5'b01111; w[5][87] = 5'b00000; w[5][88] = 5'b01111; w[5][89] = 5'b01111; w[5][90] = 5'b10000; w[5][91] = 5'b10000; w[5][92] = 5'b01111; w[5][93] = 5'b01111; w[5][94] = 5'b01111; w[5][95] = 5'b01111; w[5][96] = 5'b01111; w[5][97] = 5'b01111; w[5][98] = 5'b01111; w[5][99] = 5'b01111; w[5][100] = 5'b01111; w[5][101] = 5'b00000; w[5][102] = 5'b01111; w[5][103] = 5'b01111; w[5][104] = 5'b10000; w[5][105] = 5'b10000; w[5][106] = 5'b01111; w[5][107] = 5'b00000; w[5][108] = 5'b00000; w[5][109] = 5'b01111; w[5][110] = 5'b01111; w[5][111] = 5'b01111; w[5][112] = 5'b01111; w[5][113] = 5'b01111; w[5][114] = 5'b01111; w[5][115] = 5'b00000; w[5][116] = 5'b01111; w[5][117] = 5'b01111; w[5][118] = 5'b10000; w[5][119] = 5'b10000; w[5][120] = 5'b00000; w[5][121] = 5'b00000; w[5][122] = 5'b00000; w[5][123] = 5'b01111; w[5][124] = 5'b01111; w[5][125] = 5'b01111; w[5][126] = 5'b01111; w[5][127] = 5'b01111; w[5][128] = 5'b01111; w[5][129] = 5'b00000; w[5][130] = 5'b01111; w[5][131] = 5'b01111; w[5][132] = 5'b00000; w[5][133] = 5'b10000; w[5][134] = 5'b01111; w[5][135] = 5'b01111; w[5][136] = 5'b00000; w[5][137] = 5'b01111; w[5][138] = 5'b01111; w[5][139] = 5'b01111; w[5][140] = 5'b01111; w[5][141] = 5'b01111; w[5][142] = 5'b01111; w[5][143] = 5'b00000; w[5][144] = 5'b00000; w[5][145] = 5'b01111; w[5][146] = 5'b00000; w[5][147] = 5'b10000; w[5][148] = 5'b01111; w[5][149] = 5'b00000; w[5][150] = 5'b00000; w[5][151] = 5'b01111; w[5][152] = 5'b01111; w[5][153] = 5'b01111; w[5][154] = 5'b01111; w[5][155] = 5'b01111; w[5][156] = 5'b01111; w[5][157] = 5'b00000; w[5][158] = 5'b00000; w[5][159] = 5'b00000; w[5][160] = 5'b10000; w[5][161] = 5'b10000; w[5][162] = 5'b10000; w[5][163] = 5'b00000; w[5][164] = 5'b00000; w[5][165] = 5'b01111; w[5][166] = 5'b01111; w[5][167] = 5'b01111; w[5][168] = 5'b01111; w[5][169] = 5'b01111; w[5][170] = 5'b01111; w[5][171] = 5'b01111; w[5][172] = 5'b00000; w[5][173] = 5'b00000; w[5][174] = 5'b10000; w[5][175] = 5'b10000; w[5][176] = 5'b10000; w[5][177] = 5'b00000; w[5][178] = 5'b01111; w[5][179] = 5'b01111; w[5][180] = 5'b01111; w[5][181] = 5'b01111; w[5][182] = 5'b01111; w[5][183] = 5'b01111; w[5][184] = 5'b01111; w[5][185] = 5'b01111; w[5][186] = 5'b01111; w[5][187] = 5'b01111; w[5][188] = 5'b01111; w[5][189] = 5'b01111; w[5][190] = 5'b01111; w[5][191] = 5'b01111; w[5][192] = 5'b01111; w[5][193] = 5'b01111; w[5][194] = 5'b01111; w[5][195] = 5'b01111; w[5][196] = 5'b01111; w[5][197] = 5'b01111; w[5][198] = 5'b01111; w[5][199] = 5'b01111; w[5][200] = 5'b01111; w[5][201] = 5'b01111; w[5][202] = 5'b01111; w[5][203] = 5'b01111; w[5][204] = 5'b01111; w[5][205] = 5'b01111; w[5][206] = 5'b01111; w[5][207] = 5'b01111; w[5][208] = 5'b01111; w[5][209] = 5'b01111; 
w[6][0] = 5'b01111; w[6][1] = 5'b01111; w[6][2] = 5'b01111; w[6][3] = 5'b01111; w[6][4] = 5'b01111; w[6][5] = 5'b01111; w[6][6] = 5'b00000; w[6][7] = 5'b01111; w[6][8] = 5'b01111; w[6][9] = 5'b01111; w[6][10] = 5'b01111; w[6][11] = 5'b01111; w[6][12] = 5'b01111; w[6][13] = 5'b01111; w[6][14] = 5'b01111; w[6][15] = 5'b01111; w[6][16] = 5'b01111; w[6][17] = 5'b01111; w[6][18] = 5'b01111; w[6][19] = 5'b01111; w[6][20] = 5'b01111; w[6][21] = 5'b01111; w[6][22] = 5'b01111; w[6][23] = 5'b01111; w[6][24] = 5'b01111; w[6][25] = 5'b01111; w[6][26] = 5'b01111; w[6][27] = 5'b01111; w[6][28] = 5'b01111; w[6][29] = 5'b01111; w[6][30] = 5'b01111; w[6][31] = 5'b00000; w[6][32] = 5'b10000; w[6][33] = 5'b10000; w[6][34] = 5'b10000; w[6][35] = 5'b10000; w[6][36] = 5'b10000; w[6][37] = 5'b10000; w[6][38] = 5'b00000; w[6][39] = 5'b01111; w[6][40] = 5'b01111; w[6][41] = 5'b01111; w[6][42] = 5'b01111; w[6][43] = 5'b01111; w[6][44] = 5'b01111; w[6][45] = 5'b10000; w[6][46] = 5'b10000; w[6][47] = 5'b10000; w[6][48] = 5'b10000; w[6][49] = 5'b10000; w[6][50] = 5'b10000; w[6][51] = 5'b10000; w[6][52] = 5'b10000; w[6][53] = 5'b01111; w[6][54] = 5'b01111; w[6][55] = 5'b01111; w[6][56] = 5'b01111; w[6][57] = 5'b01111; w[6][58] = 5'b01111; w[6][59] = 5'b00000; w[6][60] = 5'b00000; w[6][61] = 5'b01111; w[6][62] = 5'b10000; w[6][63] = 5'b00000; w[6][64] = 5'b01111; w[6][65] = 5'b00000; w[6][66] = 5'b00000; w[6][67] = 5'b01111; w[6][68] = 5'b01111; w[6][69] = 5'b01111; w[6][70] = 5'b01111; w[6][71] = 5'b01111; w[6][72] = 5'b01111; w[6][73] = 5'b00000; w[6][74] = 5'b01111; w[6][75] = 5'b01111; w[6][76] = 5'b10000; w[6][77] = 5'b00000; w[6][78] = 5'b01111; w[6][79] = 5'b01111; w[6][80] = 5'b00000; w[6][81] = 5'b01111; w[6][82] = 5'b01111; w[6][83] = 5'b01111; w[6][84] = 5'b01111; w[6][85] = 5'b01111; w[6][86] = 5'b01111; w[6][87] = 5'b00000; w[6][88] = 5'b01111; w[6][89] = 5'b01111; w[6][90] = 5'b10000; w[6][91] = 5'b10000; w[6][92] = 5'b01111; w[6][93] = 5'b01111; w[6][94] = 5'b01111; w[6][95] = 5'b01111; w[6][96] = 5'b01111; w[6][97] = 5'b01111; w[6][98] = 5'b01111; w[6][99] = 5'b01111; w[6][100] = 5'b01111; w[6][101] = 5'b00000; w[6][102] = 5'b01111; w[6][103] = 5'b01111; w[6][104] = 5'b10000; w[6][105] = 5'b10000; w[6][106] = 5'b01111; w[6][107] = 5'b00000; w[6][108] = 5'b00000; w[6][109] = 5'b01111; w[6][110] = 5'b01111; w[6][111] = 5'b01111; w[6][112] = 5'b01111; w[6][113] = 5'b01111; w[6][114] = 5'b01111; w[6][115] = 5'b00000; w[6][116] = 5'b01111; w[6][117] = 5'b01111; w[6][118] = 5'b10000; w[6][119] = 5'b10000; w[6][120] = 5'b00000; w[6][121] = 5'b00000; w[6][122] = 5'b00000; w[6][123] = 5'b01111; w[6][124] = 5'b01111; w[6][125] = 5'b01111; w[6][126] = 5'b01111; w[6][127] = 5'b01111; w[6][128] = 5'b01111; w[6][129] = 5'b00000; w[6][130] = 5'b01111; w[6][131] = 5'b01111; w[6][132] = 5'b00000; w[6][133] = 5'b10000; w[6][134] = 5'b01111; w[6][135] = 5'b01111; w[6][136] = 5'b00000; w[6][137] = 5'b01111; w[6][138] = 5'b01111; w[6][139] = 5'b01111; w[6][140] = 5'b01111; w[6][141] = 5'b01111; w[6][142] = 5'b01111; w[6][143] = 5'b00000; w[6][144] = 5'b00000; w[6][145] = 5'b01111; w[6][146] = 5'b00000; w[6][147] = 5'b10000; w[6][148] = 5'b01111; w[6][149] = 5'b00000; w[6][150] = 5'b00000; w[6][151] = 5'b01111; w[6][152] = 5'b01111; w[6][153] = 5'b01111; w[6][154] = 5'b01111; w[6][155] = 5'b01111; w[6][156] = 5'b01111; w[6][157] = 5'b00000; w[6][158] = 5'b00000; w[6][159] = 5'b00000; w[6][160] = 5'b10000; w[6][161] = 5'b10000; w[6][162] = 5'b10000; w[6][163] = 5'b00000; w[6][164] = 5'b00000; w[6][165] = 5'b01111; w[6][166] = 5'b01111; w[6][167] = 5'b01111; w[6][168] = 5'b01111; w[6][169] = 5'b01111; w[6][170] = 5'b01111; w[6][171] = 5'b01111; w[6][172] = 5'b00000; w[6][173] = 5'b00000; w[6][174] = 5'b10000; w[6][175] = 5'b10000; w[6][176] = 5'b10000; w[6][177] = 5'b00000; w[6][178] = 5'b01111; w[6][179] = 5'b01111; w[6][180] = 5'b01111; w[6][181] = 5'b01111; w[6][182] = 5'b01111; w[6][183] = 5'b01111; w[6][184] = 5'b01111; w[6][185] = 5'b01111; w[6][186] = 5'b01111; w[6][187] = 5'b01111; w[6][188] = 5'b01111; w[6][189] = 5'b01111; w[6][190] = 5'b01111; w[6][191] = 5'b01111; w[6][192] = 5'b01111; w[6][193] = 5'b01111; w[6][194] = 5'b01111; w[6][195] = 5'b01111; w[6][196] = 5'b01111; w[6][197] = 5'b01111; w[6][198] = 5'b01111; w[6][199] = 5'b01111; w[6][200] = 5'b01111; w[6][201] = 5'b01111; w[6][202] = 5'b01111; w[6][203] = 5'b01111; w[6][204] = 5'b01111; w[6][205] = 5'b01111; w[6][206] = 5'b01111; w[6][207] = 5'b01111; w[6][208] = 5'b01111; w[6][209] = 5'b01111; 
w[7][0] = 5'b01111; w[7][1] = 5'b01111; w[7][2] = 5'b01111; w[7][3] = 5'b01111; w[7][4] = 5'b01111; w[7][5] = 5'b01111; w[7][6] = 5'b01111; w[7][7] = 5'b00000; w[7][8] = 5'b01111; w[7][9] = 5'b01111; w[7][10] = 5'b01111; w[7][11] = 5'b01111; w[7][12] = 5'b01111; w[7][13] = 5'b01111; w[7][14] = 5'b01111; w[7][15] = 5'b01111; w[7][16] = 5'b01111; w[7][17] = 5'b01111; w[7][18] = 5'b01111; w[7][19] = 5'b01111; w[7][20] = 5'b01111; w[7][21] = 5'b01111; w[7][22] = 5'b01111; w[7][23] = 5'b01111; w[7][24] = 5'b01111; w[7][25] = 5'b01111; w[7][26] = 5'b01111; w[7][27] = 5'b01111; w[7][28] = 5'b01111; w[7][29] = 5'b01111; w[7][30] = 5'b01111; w[7][31] = 5'b00000; w[7][32] = 5'b10000; w[7][33] = 5'b10000; w[7][34] = 5'b10000; w[7][35] = 5'b10000; w[7][36] = 5'b10000; w[7][37] = 5'b10000; w[7][38] = 5'b00000; w[7][39] = 5'b01111; w[7][40] = 5'b01111; w[7][41] = 5'b01111; w[7][42] = 5'b01111; w[7][43] = 5'b01111; w[7][44] = 5'b01111; w[7][45] = 5'b10000; w[7][46] = 5'b10000; w[7][47] = 5'b10000; w[7][48] = 5'b10000; w[7][49] = 5'b10000; w[7][50] = 5'b10000; w[7][51] = 5'b10000; w[7][52] = 5'b10000; w[7][53] = 5'b01111; w[7][54] = 5'b01111; w[7][55] = 5'b01111; w[7][56] = 5'b01111; w[7][57] = 5'b01111; w[7][58] = 5'b01111; w[7][59] = 5'b00000; w[7][60] = 5'b00000; w[7][61] = 5'b01111; w[7][62] = 5'b10000; w[7][63] = 5'b00000; w[7][64] = 5'b01111; w[7][65] = 5'b00000; w[7][66] = 5'b00000; w[7][67] = 5'b01111; w[7][68] = 5'b01111; w[7][69] = 5'b01111; w[7][70] = 5'b01111; w[7][71] = 5'b01111; w[7][72] = 5'b01111; w[7][73] = 5'b00000; w[7][74] = 5'b01111; w[7][75] = 5'b01111; w[7][76] = 5'b10000; w[7][77] = 5'b00000; w[7][78] = 5'b01111; w[7][79] = 5'b01111; w[7][80] = 5'b00000; w[7][81] = 5'b01111; w[7][82] = 5'b01111; w[7][83] = 5'b01111; w[7][84] = 5'b01111; w[7][85] = 5'b01111; w[7][86] = 5'b01111; w[7][87] = 5'b00000; w[7][88] = 5'b01111; w[7][89] = 5'b01111; w[7][90] = 5'b10000; w[7][91] = 5'b10000; w[7][92] = 5'b01111; w[7][93] = 5'b01111; w[7][94] = 5'b01111; w[7][95] = 5'b01111; w[7][96] = 5'b01111; w[7][97] = 5'b01111; w[7][98] = 5'b01111; w[7][99] = 5'b01111; w[7][100] = 5'b01111; w[7][101] = 5'b00000; w[7][102] = 5'b01111; w[7][103] = 5'b01111; w[7][104] = 5'b10000; w[7][105] = 5'b10000; w[7][106] = 5'b01111; w[7][107] = 5'b00000; w[7][108] = 5'b00000; w[7][109] = 5'b01111; w[7][110] = 5'b01111; w[7][111] = 5'b01111; w[7][112] = 5'b01111; w[7][113] = 5'b01111; w[7][114] = 5'b01111; w[7][115] = 5'b00000; w[7][116] = 5'b01111; w[7][117] = 5'b01111; w[7][118] = 5'b10000; w[7][119] = 5'b10000; w[7][120] = 5'b00000; w[7][121] = 5'b00000; w[7][122] = 5'b00000; w[7][123] = 5'b01111; w[7][124] = 5'b01111; w[7][125] = 5'b01111; w[7][126] = 5'b01111; w[7][127] = 5'b01111; w[7][128] = 5'b01111; w[7][129] = 5'b00000; w[7][130] = 5'b01111; w[7][131] = 5'b01111; w[7][132] = 5'b00000; w[7][133] = 5'b10000; w[7][134] = 5'b01111; w[7][135] = 5'b01111; w[7][136] = 5'b00000; w[7][137] = 5'b01111; w[7][138] = 5'b01111; w[7][139] = 5'b01111; w[7][140] = 5'b01111; w[7][141] = 5'b01111; w[7][142] = 5'b01111; w[7][143] = 5'b00000; w[7][144] = 5'b00000; w[7][145] = 5'b01111; w[7][146] = 5'b00000; w[7][147] = 5'b10000; w[7][148] = 5'b01111; w[7][149] = 5'b00000; w[7][150] = 5'b00000; w[7][151] = 5'b01111; w[7][152] = 5'b01111; w[7][153] = 5'b01111; w[7][154] = 5'b01111; w[7][155] = 5'b01111; w[7][156] = 5'b01111; w[7][157] = 5'b00000; w[7][158] = 5'b00000; w[7][159] = 5'b00000; w[7][160] = 5'b10000; w[7][161] = 5'b10000; w[7][162] = 5'b10000; w[7][163] = 5'b00000; w[7][164] = 5'b00000; w[7][165] = 5'b01111; w[7][166] = 5'b01111; w[7][167] = 5'b01111; w[7][168] = 5'b01111; w[7][169] = 5'b01111; w[7][170] = 5'b01111; w[7][171] = 5'b01111; w[7][172] = 5'b00000; w[7][173] = 5'b00000; w[7][174] = 5'b10000; w[7][175] = 5'b10000; w[7][176] = 5'b10000; w[7][177] = 5'b00000; w[7][178] = 5'b01111; w[7][179] = 5'b01111; w[7][180] = 5'b01111; w[7][181] = 5'b01111; w[7][182] = 5'b01111; w[7][183] = 5'b01111; w[7][184] = 5'b01111; w[7][185] = 5'b01111; w[7][186] = 5'b01111; w[7][187] = 5'b01111; w[7][188] = 5'b01111; w[7][189] = 5'b01111; w[7][190] = 5'b01111; w[7][191] = 5'b01111; w[7][192] = 5'b01111; w[7][193] = 5'b01111; w[7][194] = 5'b01111; w[7][195] = 5'b01111; w[7][196] = 5'b01111; w[7][197] = 5'b01111; w[7][198] = 5'b01111; w[7][199] = 5'b01111; w[7][200] = 5'b01111; w[7][201] = 5'b01111; w[7][202] = 5'b01111; w[7][203] = 5'b01111; w[7][204] = 5'b01111; w[7][205] = 5'b01111; w[7][206] = 5'b01111; w[7][207] = 5'b01111; w[7][208] = 5'b01111; w[7][209] = 5'b01111; 
w[8][0] = 5'b01111; w[8][1] = 5'b01111; w[8][2] = 5'b01111; w[8][3] = 5'b01111; w[8][4] = 5'b01111; w[8][5] = 5'b01111; w[8][6] = 5'b01111; w[8][7] = 5'b01111; w[8][8] = 5'b00000; w[8][9] = 5'b01111; w[8][10] = 5'b01111; w[8][11] = 5'b01111; w[8][12] = 5'b01111; w[8][13] = 5'b01111; w[8][14] = 5'b01111; w[8][15] = 5'b01111; w[8][16] = 5'b01111; w[8][17] = 5'b01111; w[8][18] = 5'b01111; w[8][19] = 5'b01111; w[8][20] = 5'b01111; w[8][21] = 5'b01111; w[8][22] = 5'b01111; w[8][23] = 5'b01111; w[8][24] = 5'b01111; w[8][25] = 5'b01111; w[8][26] = 5'b01111; w[8][27] = 5'b01111; w[8][28] = 5'b01111; w[8][29] = 5'b01111; w[8][30] = 5'b01111; w[8][31] = 5'b00000; w[8][32] = 5'b10000; w[8][33] = 5'b10000; w[8][34] = 5'b10000; w[8][35] = 5'b10000; w[8][36] = 5'b10000; w[8][37] = 5'b10000; w[8][38] = 5'b00000; w[8][39] = 5'b01111; w[8][40] = 5'b01111; w[8][41] = 5'b01111; w[8][42] = 5'b01111; w[8][43] = 5'b01111; w[8][44] = 5'b01111; w[8][45] = 5'b10000; w[8][46] = 5'b10000; w[8][47] = 5'b10000; w[8][48] = 5'b10000; w[8][49] = 5'b10000; w[8][50] = 5'b10000; w[8][51] = 5'b10000; w[8][52] = 5'b10000; w[8][53] = 5'b01111; w[8][54] = 5'b01111; w[8][55] = 5'b01111; w[8][56] = 5'b01111; w[8][57] = 5'b01111; w[8][58] = 5'b01111; w[8][59] = 5'b00000; w[8][60] = 5'b00000; w[8][61] = 5'b01111; w[8][62] = 5'b10000; w[8][63] = 5'b00000; w[8][64] = 5'b01111; w[8][65] = 5'b00000; w[8][66] = 5'b00000; w[8][67] = 5'b01111; w[8][68] = 5'b01111; w[8][69] = 5'b01111; w[8][70] = 5'b01111; w[8][71] = 5'b01111; w[8][72] = 5'b01111; w[8][73] = 5'b00000; w[8][74] = 5'b01111; w[8][75] = 5'b01111; w[8][76] = 5'b10000; w[8][77] = 5'b00000; w[8][78] = 5'b01111; w[8][79] = 5'b01111; w[8][80] = 5'b00000; w[8][81] = 5'b01111; w[8][82] = 5'b01111; w[8][83] = 5'b01111; w[8][84] = 5'b01111; w[8][85] = 5'b01111; w[8][86] = 5'b01111; w[8][87] = 5'b00000; w[8][88] = 5'b01111; w[8][89] = 5'b01111; w[8][90] = 5'b10000; w[8][91] = 5'b10000; w[8][92] = 5'b01111; w[8][93] = 5'b01111; w[8][94] = 5'b01111; w[8][95] = 5'b01111; w[8][96] = 5'b01111; w[8][97] = 5'b01111; w[8][98] = 5'b01111; w[8][99] = 5'b01111; w[8][100] = 5'b01111; w[8][101] = 5'b00000; w[8][102] = 5'b01111; w[8][103] = 5'b01111; w[8][104] = 5'b10000; w[8][105] = 5'b10000; w[8][106] = 5'b01111; w[8][107] = 5'b00000; w[8][108] = 5'b00000; w[8][109] = 5'b01111; w[8][110] = 5'b01111; w[8][111] = 5'b01111; w[8][112] = 5'b01111; w[8][113] = 5'b01111; w[8][114] = 5'b01111; w[8][115] = 5'b00000; w[8][116] = 5'b01111; w[8][117] = 5'b01111; w[8][118] = 5'b10000; w[8][119] = 5'b10000; w[8][120] = 5'b00000; w[8][121] = 5'b00000; w[8][122] = 5'b00000; w[8][123] = 5'b01111; w[8][124] = 5'b01111; w[8][125] = 5'b01111; w[8][126] = 5'b01111; w[8][127] = 5'b01111; w[8][128] = 5'b01111; w[8][129] = 5'b00000; w[8][130] = 5'b01111; w[8][131] = 5'b01111; w[8][132] = 5'b00000; w[8][133] = 5'b10000; w[8][134] = 5'b01111; w[8][135] = 5'b01111; w[8][136] = 5'b00000; w[8][137] = 5'b01111; w[8][138] = 5'b01111; w[8][139] = 5'b01111; w[8][140] = 5'b01111; w[8][141] = 5'b01111; w[8][142] = 5'b01111; w[8][143] = 5'b00000; w[8][144] = 5'b00000; w[8][145] = 5'b01111; w[8][146] = 5'b00000; w[8][147] = 5'b10000; w[8][148] = 5'b01111; w[8][149] = 5'b00000; w[8][150] = 5'b00000; w[8][151] = 5'b01111; w[8][152] = 5'b01111; w[8][153] = 5'b01111; w[8][154] = 5'b01111; w[8][155] = 5'b01111; w[8][156] = 5'b01111; w[8][157] = 5'b00000; w[8][158] = 5'b00000; w[8][159] = 5'b00000; w[8][160] = 5'b10000; w[8][161] = 5'b10000; w[8][162] = 5'b10000; w[8][163] = 5'b00000; w[8][164] = 5'b00000; w[8][165] = 5'b01111; w[8][166] = 5'b01111; w[8][167] = 5'b01111; w[8][168] = 5'b01111; w[8][169] = 5'b01111; w[8][170] = 5'b01111; w[8][171] = 5'b01111; w[8][172] = 5'b00000; w[8][173] = 5'b00000; w[8][174] = 5'b10000; w[8][175] = 5'b10000; w[8][176] = 5'b10000; w[8][177] = 5'b00000; w[8][178] = 5'b01111; w[8][179] = 5'b01111; w[8][180] = 5'b01111; w[8][181] = 5'b01111; w[8][182] = 5'b01111; w[8][183] = 5'b01111; w[8][184] = 5'b01111; w[8][185] = 5'b01111; w[8][186] = 5'b01111; w[8][187] = 5'b01111; w[8][188] = 5'b01111; w[8][189] = 5'b01111; w[8][190] = 5'b01111; w[8][191] = 5'b01111; w[8][192] = 5'b01111; w[8][193] = 5'b01111; w[8][194] = 5'b01111; w[8][195] = 5'b01111; w[8][196] = 5'b01111; w[8][197] = 5'b01111; w[8][198] = 5'b01111; w[8][199] = 5'b01111; w[8][200] = 5'b01111; w[8][201] = 5'b01111; w[8][202] = 5'b01111; w[8][203] = 5'b01111; w[8][204] = 5'b01111; w[8][205] = 5'b01111; w[8][206] = 5'b01111; w[8][207] = 5'b01111; w[8][208] = 5'b01111; w[8][209] = 5'b01111; 
w[9][0] = 5'b01111; w[9][1] = 5'b01111; w[9][2] = 5'b01111; w[9][3] = 5'b01111; w[9][4] = 5'b01111; w[9][5] = 5'b01111; w[9][6] = 5'b01111; w[9][7] = 5'b01111; w[9][8] = 5'b01111; w[9][9] = 5'b00000; w[9][10] = 5'b01111; w[9][11] = 5'b01111; w[9][12] = 5'b01111; w[9][13] = 5'b01111; w[9][14] = 5'b01111; w[9][15] = 5'b01111; w[9][16] = 5'b01111; w[9][17] = 5'b01111; w[9][18] = 5'b01111; w[9][19] = 5'b01111; w[9][20] = 5'b01111; w[9][21] = 5'b01111; w[9][22] = 5'b01111; w[9][23] = 5'b01111; w[9][24] = 5'b01111; w[9][25] = 5'b01111; w[9][26] = 5'b01111; w[9][27] = 5'b01111; w[9][28] = 5'b01111; w[9][29] = 5'b01111; w[9][30] = 5'b01111; w[9][31] = 5'b00000; w[9][32] = 5'b10000; w[9][33] = 5'b10000; w[9][34] = 5'b10000; w[9][35] = 5'b10000; w[9][36] = 5'b10000; w[9][37] = 5'b10000; w[9][38] = 5'b00000; w[9][39] = 5'b01111; w[9][40] = 5'b01111; w[9][41] = 5'b01111; w[9][42] = 5'b01111; w[9][43] = 5'b01111; w[9][44] = 5'b01111; w[9][45] = 5'b10000; w[9][46] = 5'b10000; w[9][47] = 5'b10000; w[9][48] = 5'b10000; w[9][49] = 5'b10000; w[9][50] = 5'b10000; w[9][51] = 5'b10000; w[9][52] = 5'b10000; w[9][53] = 5'b01111; w[9][54] = 5'b01111; w[9][55] = 5'b01111; w[9][56] = 5'b01111; w[9][57] = 5'b01111; w[9][58] = 5'b01111; w[9][59] = 5'b00000; w[9][60] = 5'b00000; w[9][61] = 5'b01111; w[9][62] = 5'b10000; w[9][63] = 5'b00000; w[9][64] = 5'b01111; w[9][65] = 5'b00000; w[9][66] = 5'b00000; w[9][67] = 5'b01111; w[9][68] = 5'b01111; w[9][69] = 5'b01111; w[9][70] = 5'b01111; w[9][71] = 5'b01111; w[9][72] = 5'b01111; w[9][73] = 5'b00000; w[9][74] = 5'b01111; w[9][75] = 5'b01111; w[9][76] = 5'b10000; w[9][77] = 5'b00000; w[9][78] = 5'b01111; w[9][79] = 5'b01111; w[9][80] = 5'b00000; w[9][81] = 5'b01111; w[9][82] = 5'b01111; w[9][83] = 5'b01111; w[9][84] = 5'b01111; w[9][85] = 5'b01111; w[9][86] = 5'b01111; w[9][87] = 5'b00000; w[9][88] = 5'b01111; w[9][89] = 5'b01111; w[9][90] = 5'b10000; w[9][91] = 5'b10000; w[9][92] = 5'b01111; w[9][93] = 5'b01111; w[9][94] = 5'b01111; w[9][95] = 5'b01111; w[9][96] = 5'b01111; w[9][97] = 5'b01111; w[9][98] = 5'b01111; w[9][99] = 5'b01111; w[9][100] = 5'b01111; w[9][101] = 5'b00000; w[9][102] = 5'b01111; w[9][103] = 5'b01111; w[9][104] = 5'b10000; w[9][105] = 5'b10000; w[9][106] = 5'b01111; w[9][107] = 5'b00000; w[9][108] = 5'b00000; w[9][109] = 5'b01111; w[9][110] = 5'b01111; w[9][111] = 5'b01111; w[9][112] = 5'b01111; w[9][113] = 5'b01111; w[9][114] = 5'b01111; w[9][115] = 5'b00000; w[9][116] = 5'b01111; w[9][117] = 5'b01111; w[9][118] = 5'b10000; w[9][119] = 5'b10000; w[9][120] = 5'b00000; w[9][121] = 5'b00000; w[9][122] = 5'b00000; w[9][123] = 5'b01111; w[9][124] = 5'b01111; w[9][125] = 5'b01111; w[9][126] = 5'b01111; w[9][127] = 5'b01111; w[9][128] = 5'b01111; w[9][129] = 5'b00000; w[9][130] = 5'b01111; w[9][131] = 5'b01111; w[9][132] = 5'b00000; w[9][133] = 5'b10000; w[9][134] = 5'b01111; w[9][135] = 5'b01111; w[9][136] = 5'b00000; w[9][137] = 5'b01111; w[9][138] = 5'b01111; w[9][139] = 5'b01111; w[9][140] = 5'b01111; w[9][141] = 5'b01111; w[9][142] = 5'b01111; w[9][143] = 5'b00000; w[9][144] = 5'b00000; w[9][145] = 5'b01111; w[9][146] = 5'b00000; w[9][147] = 5'b10000; w[9][148] = 5'b01111; w[9][149] = 5'b00000; w[9][150] = 5'b00000; w[9][151] = 5'b01111; w[9][152] = 5'b01111; w[9][153] = 5'b01111; w[9][154] = 5'b01111; w[9][155] = 5'b01111; w[9][156] = 5'b01111; w[9][157] = 5'b00000; w[9][158] = 5'b00000; w[9][159] = 5'b00000; w[9][160] = 5'b10000; w[9][161] = 5'b10000; w[9][162] = 5'b10000; w[9][163] = 5'b00000; w[9][164] = 5'b00000; w[9][165] = 5'b01111; w[9][166] = 5'b01111; w[9][167] = 5'b01111; w[9][168] = 5'b01111; w[9][169] = 5'b01111; w[9][170] = 5'b01111; w[9][171] = 5'b01111; w[9][172] = 5'b00000; w[9][173] = 5'b00000; w[9][174] = 5'b10000; w[9][175] = 5'b10000; w[9][176] = 5'b10000; w[9][177] = 5'b00000; w[9][178] = 5'b01111; w[9][179] = 5'b01111; w[9][180] = 5'b01111; w[9][181] = 5'b01111; w[9][182] = 5'b01111; w[9][183] = 5'b01111; w[9][184] = 5'b01111; w[9][185] = 5'b01111; w[9][186] = 5'b01111; w[9][187] = 5'b01111; w[9][188] = 5'b01111; w[9][189] = 5'b01111; w[9][190] = 5'b01111; w[9][191] = 5'b01111; w[9][192] = 5'b01111; w[9][193] = 5'b01111; w[9][194] = 5'b01111; w[9][195] = 5'b01111; w[9][196] = 5'b01111; w[9][197] = 5'b01111; w[9][198] = 5'b01111; w[9][199] = 5'b01111; w[9][200] = 5'b01111; w[9][201] = 5'b01111; w[9][202] = 5'b01111; w[9][203] = 5'b01111; w[9][204] = 5'b01111; w[9][205] = 5'b01111; w[9][206] = 5'b01111; w[9][207] = 5'b01111; w[9][208] = 5'b01111; w[9][209] = 5'b01111; 
w[10][0] = 5'b01111; w[10][1] = 5'b01111; w[10][2] = 5'b01111; w[10][3] = 5'b01111; w[10][4] = 5'b01111; w[10][5] = 5'b01111; w[10][6] = 5'b01111; w[10][7] = 5'b01111; w[10][8] = 5'b01111; w[10][9] = 5'b01111; w[10][10] = 5'b00000; w[10][11] = 5'b01111; w[10][12] = 5'b01111; w[10][13] = 5'b01111; w[10][14] = 5'b01111; w[10][15] = 5'b01111; w[10][16] = 5'b01111; w[10][17] = 5'b01111; w[10][18] = 5'b01111; w[10][19] = 5'b01111; w[10][20] = 5'b01111; w[10][21] = 5'b01111; w[10][22] = 5'b01111; w[10][23] = 5'b01111; w[10][24] = 5'b01111; w[10][25] = 5'b01111; w[10][26] = 5'b01111; w[10][27] = 5'b01111; w[10][28] = 5'b01111; w[10][29] = 5'b01111; w[10][30] = 5'b01111; w[10][31] = 5'b00000; w[10][32] = 5'b10000; w[10][33] = 5'b10000; w[10][34] = 5'b10000; w[10][35] = 5'b10000; w[10][36] = 5'b10000; w[10][37] = 5'b10000; w[10][38] = 5'b00000; w[10][39] = 5'b01111; w[10][40] = 5'b01111; w[10][41] = 5'b01111; w[10][42] = 5'b01111; w[10][43] = 5'b01111; w[10][44] = 5'b01111; w[10][45] = 5'b10000; w[10][46] = 5'b10000; w[10][47] = 5'b10000; w[10][48] = 5'b10000; w[10][49] = 5'b10000; w[10][50] = 5'b10000; w[10][51] = 5'b10000; w[10][52] = 5'b10000; w[10][53] = 5'b01111; w[10][54] = 5'b01111; w[10][55] = 5'b01111; w[10][56] = 5'b01111; w[10][57] = 5'b01111; w[10][58] = 5'b01111; w[10][59] = 5'b00000; w[10][60] = 5'b00000; w[10][61] = 5'b01111; w[10][62] = 5'b10000; w[10][63] = 5'b00000; w[10][64] = 5'b01111; w[10][65] = 5'b00000; w[10][66] = 5'b00000; w[10][67] = 5'b01111; w[10][68] = 5'b01111; w[10][69] = 5'b01111; w[10][70] = 5'b01111; w[10][71] = 5'b01111; w[10][72] = 5'b01111; w[10][73] = 5'b00000; w[10][74] = 5'b01111; w[10][75] = 5'b01111; w[10][76] = 5'b10000; w[10][77] = 5'b00000; w[10][78] = 5'b01111; w[10][79] = 5'b01111; w[10][80] = 5'b00000; w[10][81] = 5'b01111; w[10][82] = 5'b01111; w[10][83] = 5'b01111; w[10][84] = 5'b01111; w[10][85] = 5'b01111; w[10][86] = 5'b01111; w[10][87] = 5'b00000; w[10][88] = 5'b01111; w[10][89] = 5'b01111; w[10][90] = 5'b10000; w[10][91] = 5'b10000; w[10][92] = 5'b01111; w[10][93] = 5'b01111; w[10][94] = 5'b01111; w[10][95] = 5'b01111; w[10][96] = 5'b01111; w[10][97] = 5'b01111; w[10][98] = 5'b01111; w[10][99] = 5'b01111; w[10][100] = 5'b01111; w[10][101] = 5'b00000; w[10][102] = 5'b01111; w[10][103] = 5'b01111; w[10][104] = 5'b10000; w[10][105] = 5'b10000; w[10][106] = 5'b01111; w[10][107] = 5'b00000; w[10][108] = 5'b00000; w[10][109] = 5'b01111; w[10][110] = 5'b01111; w[10][111] = 5'b01111; w[10][112] = 5'b01111; w[10][113] = 5'b01111; w[10][114] = 5'b01111; w[10][115] = 5'b00000; w[10][116] = 5'b01111; w[10][117] = 5'b01111; w[10][118] = 5'b10000; w[10][119] = 5'b10000; w[10][120] = 5'b00000; w[10][121] = 5'b00000; w[10][122] = 5'b00000; w[10][123] = 5'b01111; w[10][124] = 5'b01111; w[10][125] = 5'b01111; w[10][126] = 5'b01111; w[10][127] = 5'b01111; w[10][128] = 5'b01111; w[10][129] = 5'b00000; w[10][130] = 5'b01111; w[10][131] = 5'b01111; w[10][132] = 5'b00000; w[10][133] = 5'b10000; w[10][134] = 5'b01111; w[10][135] = 5'b01111; w[10][136] = 5'b00000; w[10][137] = 5'b01111; w[10][138] = 5'b01111; w[10][139] = 5'b01111; w[10][140] = 5'b01111; w[10][141] = 5'b01111; w[10][142] = 5'b01111; w[10][143] = 5'b00000; w[10][144] = 5'b00000; w[10][145] = 5'b01111; w[10][146] = 5'b00000; w[10][147] = 5'b10000; w[10][148] = 5'b01111; w[10][149] = 5'b00000; w[10][150] = 5'b00000; w[10][151] = 5'b01111; w[10][152] = 5'b01111; w[10][153] = 5'b01111; w[10][154] = 5'b01111; w[10][155] = 5'b01111; w[10][156] = 5'b01111; w[10][157] = 5'b00000; w[10][158] = 5'b00000; w[10][159] = 5'b00000; w[10][160] = 5'b10000; w[10][161] = 5'b10000; w[10][162] = 5'b10000; w[10][163] = 5'b00000; w[10][164] = 5'b00000; w[10][165] = 5'b01111; w[10][166] = 5'b01111; w[10][167] = 5'b01111; w[10][168] = 5'b01111; w[10][169] = 5'b01111; w[10][170] = 5'b01111; w[10][171] = 5'b01111; w[10][172] = 5'b00000; w[10][173] = 5'b00000; w[10][174] = 5'b10000; w[10][175] = 5'b10000; w[10][176] = 5'b10000; w[10][177] = 5'b00000; w[10][178] = 5'b01111; w[10][179] = 5'b01111; w[10][180] = 5'b01111; w[10][181] = 5'b01111; w[10][182] = 5'b01111; w[10][183] = 5'b01111; w[10][184] = 5'b01111; w[10][185] = 5'b01111; w[10][186] = 5'b01111; w[10][187] = 5'b01111; w[10][188] = 5'b01111; w[10][189] = 5'b01111; w[10][190] = 5'b01111; w[10][191] = 5'b01111; w[10][192] = 5'b01111; w[10][193] = 5'b01111; w[10][194] = 5'b01111; w[10][195] = 5'b01111; w[10][196] = 5'b01111; w[10][197] = 5'b01111; w[10][198] = 5'b01111; w[10][199] = 5'b01111; w[10][200] = 5'b01111; w[10][201] = 5'b01111; w[10][202] = 5'b01111; w[10][203] = 5'b01111; w[10][204] = 5'b01111; w[10][205] = 5'b01111; w[10][206] = 5'b01111; w[10][207] = 5'b01111; w[10][208] = 5'b01111; w[10][209] = 5'b01111; 
w[11][0] = 5'b01111; w[11][1] = 5'b01111; w[11][2] = 5'b01111; w[11][3] = 5'b01111; w[11][4] = 5'b01111; w[11][5] = 5'b01111; w[11][6] = 5'b01111; w[11][7] = 5'b01111; w[11][8] = 5'b01111; w[11][9] = 5'b01111; w[11][10] = 5'b01111; w[11][11] = 5'b00000; w[11][12] = 5'b01111; w[11][13] = 5'b01111; w[11][14] = 5'b01111; w[11][15] = 5'b01111; w[11][16] = 5'b01111; w[11][17] = 5'b01111; w[11][18] = 5'b01111; w[11][19] = 5'b01111; w[11][20] = 5'b01111; w[11][21] = 5'b01111; w[11][22] = 5'b01111; w[11][23] = 5'b01111; w[11][24] = 5'b01111; w[11][25] = 5'b01111; w[11][26] = 5'b01111; w[11][27] = 5'b01111; w[11][28] = 5'b01111; w[11][29] = 5'b01111; w[11][30] = 5'b01111; w[11][31] = 5'b00000; w[11][32] = 5'b10000; w[11][33] = 5'b10000; w[11][34] = 5'b10000; w[11][35] = 5'b10000; w[11][36] = 5'b10000; w[11][37] = 5'b10000; w[11][38] = 5'b00000; w[11][39] = 5'b01111; w[11][40] = 5'b01111; w[11][41] = 5'b01111; w[11][42] = 5'b01111; w[11][43] = 5'b01111; w[11][44] = 5'b01111; w[11][45] = 5'b10000; w[11][46] = 5'b10000; w[11][47] = 5'b10000; w[11][48] = 5'b10000; w[11][49] = 5'b10000; w[11][50] = 5'b10000; w[11][51] = 5'b10000; w[11][52] = 5'b10000; w[11][53] = 5'b01111; w[11][54] = 5'b01111; w[11][55] = 5'b01111; w[11][56] = 5'b01111; w[11][57] = 5'b01111; w[11][58] = 5'b01111; w[11][59] = 5'b00000; w[11][60] = 5'b00000; w[11][61] = 5'b01111; w[11][62] = 5'b10000; w[11][63] = 5'b00000; w[11][64] = 5'b01111; w[11][65] = 5'b00000; w[11][66] = 5'b00000; w[11][67] = 5'b01111; w[11][68] = 5'b01111; w[11][69] = 5'b01111; w[11][70] = 5'b01111; w[11][71] = 5'b01111; w[11][72] = 5'b01111; w[11][73] = 5'b00000; w[11][74] = 5'b01111; w[11][75] = 5'b01111; w[11][76] = 5'b10000; w[11][77] = 5'b00000; w[11][78] = 5'b01111; w[11][79] = 5'b01111; w[11][80] = 5'b00000; w[11][81] = 5'b01111; w[11][82] = 5'b01111; w[11][83] = 5'b01111; w[11][84] = 5'b01111; w[11][85] = 5'b01111; w[11][86] = 5'b01111; w[11][87] = 5'b00000; w[11][88] = 5'b01111; w[11][89] = 5'b01111; w[11][90] = 5'b10000; w[11][91] = 5'b10000; w[11][92] = 5'b01111; w[11][93] = 5'b01111; w[11][94] = 5'b01111; w[11][95] = 5'b01111; w[11][96] = 5'b01111; w[11][97] = 5'b01111; w[11][98] = 5'b01111; w[11][99] = 5'b01111; w[11][100] = 5'b01111; w[11][101] = 5'b00000; w[11][102] = 5'b01111; w[11][103] = 5'b01111; w[11][104] = 5'b10000; w[11][105] = 5'b10000; w[11][106] = 5'b01111; w[11][107] = 5'b00000; w[11][108] = 5'b00000; w[11][109] = 5'b01111; w[11][110] = 5'b01111; w[11][111] = 5'b01111; w[11][112] = 5'b01111; w[11][113] = 5'b01111; w[11][114] = 5'b01111; w[11][115] = 5'b00000; w[11][116] = 5'b01111; w[11][117] = 5'b01111; w[11][118] = 5'b10000; w[11][119] = 5'b10000; w[11][120] = 5'b00000; w[11][121] = 5'b00000; w[11][122] = 5'b00000; w[11][123] = 5'b01111; w[11][124] = 5'b01111; w[11][125] = 5'b01111; w[11][126] = 5'b01111; w[11][127] = 5'b01111; w[11][128] = 5'b01111; w[11][129] = 5'b00000; w[11][130] = 5'b01111; w[11][131] = 5'b01111; w[11][132] = 5'b00000; w[11][133] = 5'b10000; w[11][134] = 5'b01111; w[11][135] = 5'b01111; w[11][136] = 5'b00000; w[11][137] = 5'b01111; w[11][138] = 5'b01111; w[11][139] = 5'b01111; w[11][140] = 5'b01111; w[11][141] = 5'b01111; w[11][142] = 5'b01111; w[11][143] = 5'b00000; w[11][144] = 5'b00000; w[11][145] = 5'b01111; w[11][146] = 5'b00000; w[11][147] = 5'b10000; w[11][148] = 5'b01111; w[11][149] = 5'b00000; w[11][150] = 5'b00000; w[11][151] = 5'b01111; w[11][152] = 5'b01111; w[11][153] = 5'b01111; w[11][154] = 5'b01111; w[11][155] = 5'b01111; w[11][156] = 5'b01111; w[11][157] = 5'b00000; w[11][158] = 5'b00000; w[11][159] = 5'b00000; w[11][160] = 5'b10000; w[11][161] = 5'b10000; w[11][162] = 5'b10000; w[11][163] = 5'b00000; w[11][164] = 5'b00000; w[11][165] = 5'b01111; w[11][166] = 5'b01111; w[11][167] = 5'b01111; w[11][168] = 5'b01111; w[11][169] = 5'b01111; w[11][170] = 5'b01111; w[11][171] = 5'b01111; w[11][172] = 5'b00000; w[11][173] = 5'b00000; w[11][174] = 5'b10000; w[11][175] = 5'b10000; w[11][176] = 5'b10000; w[11][177] = 5'b00000; w[11][178] = 5'b01111; w[11][179] = 5'b01111; w[11][180] = 5'b01111; w[11][181] = 5'b01111; w[11][182] = 5'b01111; w[11][183] = 5'b01111; w[11][184] = 5'b01111; w[11][185] = 5'b01111; w[11][186] = 5'b01111; w[11][187] = 5'b01111; w[11][188] = 5'b01111; w[11][189] = 5'b01111; w[11][190] = 5'b01111; w[11][191] = 5'b01111; w[11][192] = 5'b01111; w[11][193] = 5'b01111; w[11][194] = 5'b01111; w[11][195] = 5'b01111; w[11][196] = 5'b01111; w[11][197] = 5'b01111; w[11][198] = 5'b01111; w[11][199] = 5'b01111; w[11][200] = 5'b01111; w[11][201] = 5'b01111; w[11][202] = 5'b01111; w[11][203] = 5'b01111; w[11][204] = 5'b01111; w[11][205] = 5'b01111; w[11][206] = 5'b01111; w[11][207] = 5'b01111; w[11][208] = 5'b01111; w[11][209] = 5'b01111; 
w[12][0] = 5'b01111; w[12][1] = 5'b01111; w[12][2] = 5'b01111; w[12][3] = 5'b01111; w[12][4] = 5'b01111; w[12][5] = 5'b01111; w[12][6] = 5'b01111; w[12][7] = 5'b01111; w[12][8] = 5'b01111; w[12][9] = 5'b01111; w[12][10] = 5'b01111; w[12][11] = 5'b01111; w[12][12] = 5'b00000; w[12][13] = 5'b01111; w[12][14] = 5'b01111; w[12][15] = 5'b01111; w[12][16] = 5'b01111; w[12][17] = 5'b01111; w[12][18] = 5'b01111; w[12][19] = 5'b01111; w[12][20] = 5'b01111; w[12][21] = 5'b01111; w[12][22] = 5'b01111; w[12][23] = 5'b01111; w[12][24] = 5'b01111; w[12][25] = 5'b01111; w[12][26] = 5'b01111; w[12][27] = 5'b01111; w[12][28] = 5'b01111; w[12][29] = 5'b01111; w[12][30] = 5'b01111; w[12][31] = 5'b00000; w[12][32] = 5'b10000; w[12][33] = 5'b10000; w[12][34] = 5'b10000; w[12][35] = 5'b10000; w[12][36] = 5'b10000; w[12][37] = 5'b10000; w[12][38] = 5'b00000; w[12][39] = 5'b01111; w[12][40] = 5'b01111; w[12][41] = 5'b01111; w[12][42] = 5'b01111; w[12][43] = 5'b01111; w[12][44] = 5'b01111; w[12][45] = 5'b10000; w[12][46] = 5'b10000; w[12][47] = 5'b10000; w[12][48] = 5'b10000; w[12][49] = 5'b10000; w[12][50] = 5'b10000; w[12][51] = 5'b10000; w[12][52] = 5'b10000; w[12][53] = 5'b01111; w[12][54] = 5'b01111; w[12][55] = 5'b01111; w[12][56] = 5'b01111; w[12][57] = 5'b01111; w[12][58] = 5'b01111; w[12][59] = 5'b00000; w[12][60] = 5'b00000; w[12][61] = 5'b01111; w[12][62] = 5'b10000; w[12][63] = 5'b00000; w[12][64] = 5'b01111; w[12][65] = 5'b00000; w[12][66] = 5'b00000; w[12][67] = 5'b01111; w[12][68] = 5'b01111; w[12][69] = 5'b01111; w[12][70] = 5'b01111; w[12][71] = 5'b01111; w[12][72] = 5'b01111; w[12][73] = 5'b00000; w[12][74] = 5'b01111; w[12][75] = 5'b01111; w[12][76] = 5'b10000; w[12][77] = 5'b00000; w[12][78] = 5'b01111; w[12][79] = 5'b01111; w[12][80] = 5'b00000; w[12][81] = 5'b01111; w[12][82] = 5'b01111; w[12][83] = 5'b01111; w[12][84] = 5'b01111; w[12][85] = 5'b01111; w[12][86] = 5'b01111; w[12][87] = 5'b00000; w[12][88] = 5'b01111; w[12][89] = 5'b01111; w[12][90] = 5'b10000; w[12][91] = 5'b10000; w[12][92] = 5'b01111; w[12][93] = 5'b01111; w[12][94] = 5'b01111; w[12][95] = 5'b01111; w[12][96] = 5'b01111; w[12][97] = 5'b01111; w[12][98] = 5'b01111; w[12][99] = 5'b01111; w[12][100] = 5'b01111; w[12][101] = 5'b00000; w[12][102] = 5'b01111; w[12][103] = 5'b01111; w[12][104] = 5'b10000; w[12][105] = 5'b10000; w[12][106] = 5'b01111; w[12][107] = 5'b00000; w[12][108] = 5'b00000; w[12][109] = 5'b01111; w[12][110] = 5'b01111; w[12][111] = 5'b01111; w[12][112] = 5'b01111; w[12][113] = 5'b01111; w[12][114] = 5'b01111; w[12][115] = 5'b00000; w[12][116] = 5'b01111; w[12][117] = 5'b01111; w[12][118] = 5'b10000; w[12][119] = 5'b10000; w[12][120] = 5'b00000; w[12][121] = 5'b00000; w[12][122] = 5'b00000; w[12][123] = 5'b01111; w[12][124] = 5'b01111; w[12][125] = 5'b01111; w[12][126] = 5'b01111; w[12][127] = 5'b01111; w[12][128] = 5'b01111; w[12][129] = 5'b00000; w[12][130] = 5'b01111; w[12][131] = 5'b01111; w[12][132] = 5'b00000; w[12][133] = 5'b10000; w[12][134] = 5'b01111; w[12][135] = 5'b01111; w[12][136] = 5'b00000; w[12][137] = 5'b01111; w[12][138] = 5'b01111; w[12][139] = 5'b01111; w[12][140] = 5'b01111; w[12][141] = 5'b01111; w[12][142] = 5'b01111; w[12][143] = 5'b00000; w[12][144] = 5'b00000; w[12][145] = 5'b01111; w[12][146] = 5'b00000; w[12][147] = 5'b10000; w[12][148] = 5'b01111; w[12][149] = 5'b00000; w[12][150] = 5'b00000; w[12][151] = 5'b01111; w[12][152] = 5'b01111; w[12][153] = 5'b01111; w[12][154] = 5'b01111; w[12][155] = 5'b01111; w[12][156] = 5'b01111; w[12][157] = 5'b00000; w[12][158] = 5'b00000; w[12][159] = 5'b00000; w[12][160] = 5'b10000; w[12][161] = 5'b10000; w[12][162] = 5'b10000; w[12][163] = 5'b00000; w[12][164] = 5'b00000; w[12][165] = 5'b01111; w[12][166] = 5'b01111; w[12][167] = 5'b01111; w[12][168] = 5'b01111; w[12][169] = 5'b01111; w[12][170] = 5'b01111; w[12][171] = 5'b01111; w[12][172] = 5'b00000; w[12][173] = 5'b00000; w[12][174] = 5'b10000; w[12][175] = 5'b10000; w[12][176] = 5'b10000; w[12][177] = 5'b00000; w[12][178] = 5'b01111; w[12][179] = 5'b01111; w[12][180] = 5'b01111; w[12][181] = 5'b01111; w[12][182] = 5'b01111; w[12][183] = 5'b01111; w[12][184] = 5'b01111; w[12][185] = 5'b01111; w[12][186] = 5'b01111; w[12][187] = 5'b01111; w[12][188] = 5'b01111; w[12][189] = 5'b01111; w[12][190] = 5'b01111; w[12][191] = 5'b01111; w[12][192] = 5'b01111; w[12][193] = 5'b01111; w[12][194] = 5'b01111; w[12][195] = 5'b01111; w[12][196] = 5'b01111; w[12][197] = 5'b01111; w[12][198] = 5'b01111; w[12][199] = 5'b01111; w[12][200] = 5'b01111; w[12][201] = 5'b01111; w[12][202] = 5'b01111; w[12][203] = 5'b01111; w[12][204] = 5'b01111; w[12][205] = 5'b01111; w[12][206] = 5'b01111; w[12][207] = 5'b01111; w[12][208] = 5'b01111; w[12][209] = 5'b01111; 
w[13][0] = 5'b01111; w[13][1] = 5'b01111; w[13][2] = 5'b01111; w[13][3] = 5'b01111; w[13][4] = 5'b01111; w[13][5] = 5'b01111; w[13][6] = 5'b01111; w[13][7] = 5'b01111; w[13][8] = 5'b01111; w[13][9] = 5'b01111; w[13][10] = 5'b01111; w[13][11] = 5'b01111; w[13][12] = 5'b01111; w[13][13] = 5'b00000; w[13][14] = 5'b01111; w[13][15] = 5'b01111; w[13][16] = 5'b01111; w[13][17] = 5'b01111; w[13][18] = 5'b01111; w[13][19] = 5'b01111; w[13][20] = 5'b01111; w[13][21] = 5'b01111; w[13][22] = 5'b01111; w[13][23] = 5'b01111; w[13][24] = 5'b01111; w[13][25] = 5'b01111; w[13][26] = 5'b01111; w[13][27] = 5'b01111; w[13][28] = 5'b01111; w[13][29] = 5'b01111; w[13][30] = 5'b01111; w[13][31] = 5'b00000; w[13][32] = 5'b10000; w[13][33] = 5'b10000; w[13][34] = 5'b10000; w[13][35] = 5'b10000; w[13][36] = 5'b10000; w[13][37] = 5'b10000; w[13][38] = 5'b00000; w[13][39] = 5'b01111; w[13][40] = 5'b01111; w[13][41] = 5'b01111; w[13][42] = 5'b01111; w[13][43] = 5'b01111; w[13][44] = 5'b01111; w[13][45] = 5'b10000; w[13][46] = 5'b10000; w[13][47] = 5'b10000; w[13][48] = 5'b10000; w[13][49] = 5'b10000; w[13][50] = 5'b10000; w[13][51] = 5'b10000; w[13][52] = 5'b10000; w[13][53] = 5'b01111; w[13][54] = 5'b01111; w[13][55] = 5'b01111; w[13][56] = 5'b01111; w[13][57] = 5'b01111; w[13][58] = 5'b01111; w[13][59] = 5'b00000; w[13][60] = 5'b00000; w[13][61] = 5'b01111; w[13][62] = 5'b10000; w[13][63] = 5'b00000; w[13][64] = 5'b01111; w[13][65] = 5'b00000; w[13][66] = 5'b00000; w[13][67] = 5'b01111; w[13][68] = 5'b01111; w[13][69] = 5'b01111; w[13][70] = 5'b01111; w[13][71] = 5'b01111; w[13][72] = 5'b01111; w[13][73] = 5'b00000; w[13][74] = 5'b01111; w[13][75] = 5'b01111; w[13][76] = 5'b10000; w[13][77] = 5'b00000; w[13][78] = 5'b01111; w[13][79] = 5'b01111; w[13][80] = 5'b00000; w[13][81] = 5'b01111; w[13][82] = 5'b01111; w[13][83] = 5'b01111; w[13][84] = 5'b01111; w[13][85] = 5'b01111; w[13][86] = 5'b01111; w[13][87] = 5'b00000; w[13][88] = 5'b01111; w[13][89] = 5'b01111; w[13][90] = 5'b10000; w[13][91] = 5'b10000; w[13][92] = 5'b01111; w[13][93] = 5'b01111; w[13][94] = 5'b01111; w[13][95] = 5'b01111; w[13][96] = 5'b01111; w[13][97] = 5'b01111; w[13][98] = 5'b01111; w[13][99] = 5'b01111; w[13][100] = 5'b01111; w[13][101] = 5'b00000; w[13][102] = 5'b01111; w[13][103] = 5'b01111; w[13][104] = 5'b10000; w[13][105] = 5'b10000; w[13][106] = 5'b01111; w[13][107] = 5'b00000; w[13][108] = 5'b00000; w[13][109] = 5'b01111; w[13][110] = 5'b01111; w[13][111] = 5'b01111; w[13][112] = 5'b01111; w[13][113] = 5'b01111; w[13][114] = 5'b01111; w[13][115] = 5'b00000; w[13][116] = 5'b01111; w[13][117] = 5'b01111; w[13][118] = 5'b10000; w[13][119] = 5'b10000; w[13][120] = 5'b00000; w[13][121] = 5'b00000; w[13][122] = 5'b00000; w[13][123] = 5'b01111; w[13][124] = 5'b01111; w[13][125] = 5'b01111; w[13][126] = 5'b01111; w[13][127] = 5'b01111; w[13][128] = 5'b01111; w[13][129] = 5'b00000; w[13][130] = 5'b01111; w[13][131] = 5'b01111; w[13][132] = 5'b00000; w[13][133] = 5'b10000; w[13][134] = 5'b01111; w[13][135] = 5'b01111; w[13][136] = 5'b00000; w[13][137] = 5'b01111; w[13][138] = 5'b01111; w[13][139] = 5'b01111; w[13][140] = 5'b01111; w[13][141] = 5'b01111; w[13][142] = 5'b01111; w[13][143] = 5'b00000; w[13][144] = 5'b00000; w[13][145] = 5'b01111; w[13][146] = 5'b00000; w[13][147] = 5'b10000; w[13][148] = 5'b01111; w[13][149] = 5'b00000; w[13][150] = 5'b00000; w[13][151] = 5'b01111; w[13][152] = 5'b01111; w[13][153] = 5'b01111; w[13][154] = 5'b01111; w[13][155] = 5'b01111; w[13][156] = 5'b01111; w[13][157] = 5'b00000; w[13][158] = 5'b00000; w[13][159] = 5'b00000; w[13][160] = 5'b10000; w[13][161] = 5'b10000; w[13][162] = 5'b10000; w[13][163] = 5'b00000; w[13][164] = 5'b00000; w[13][165] = 5'b01111; w[13][166] = 5'b01111; w[13][167] = 5'b01111; w[13][168] = 5'b01111; w[13][169] = 5'b01111; w[13][170] = 5'b01111; w[13][171] = 5'b01111; w[13][172] = 5'b00000; w[13][173] = 5'b00000; w[13][174] = 5'b10000; w[13][175] = 5'b10000; w[13][176] = 5'b10000; w[13][177] = 5'b00000; w[13][178] = 5'b01111; w[13][179] = 5'b01111; w[13][180] = 5'b01111; w[13][181] = 5'b01111; w[13][182] = 5'b01111; w[13][183] = 5'b01111; w[13][184] = 5'b01111; w[13][185] = 5'b01111; w[13][186] = 5'b01111; w[13][187] = 5'b01111; w[13][188] = 5'b01111; w[13][189] = 5'b01111; w[13][190] = 5'b01111; w[13][191] = 5'b01111; w[13][192] = 5'b01111; w[13][193] = 5'b01111; w[13][194] = 5'b01111; w[13][195] = 5'b01111; w[13][196] = 5'b01111; w[13][197] = 5'b01111; w[13][198] = 5'b01111; w[13][199] = 5'b01111; w[13][200] = 5'b01111; w[13][201] = 5'b01111; w[13][202] = 5'b01111; w[13][203] = 5'b01111; w[13][204] = 5'b01111; w[13][205] = 5'b01111; w[13][206] = 5'b01111; w[13][207] = 5'b01111; w[13][208] = 5'b01111; w[13][209] = 5'b01111; 
w[14][0] = 5'b01111; w[14][1] = 5'b01111; w[14][2] = 5'b01111; w[14][3] = 5'b01111; w[14][4] = 5'b01111; w[14][5] = 5'b01111; w[14][6] = 5'b01111; w[14][7] = 5'b01111; w[14][8] = 5'b01111; w[14][9] = 5'b01111; w[14][10] = 5'b01111; w[14][11] = 5'b01111; w[14][12] = 5'b01111; w[14][13] = 5'b01111; w[14][14] = 5'b00000; w[14][15] = 5'b01111; w[14][16] = 5'b01111; w[14][17] = 5'b01111; w[14][18] = 5'b01111; w[14][19] = 5'b01111; w[14][20] = 5'b01111; w[14][21] = 5'b01111; w[14][22] = 5'b01111; w[14][23] = 5'b01111; w[14][24] = 5'b01111; w[14][25] = 5'b01111; w[14][26] = 5'b01111; w[14][27] = 5'b01111; w[14][28] = 5'b01111; w[14][29] = 5'b01111; w[14][30] = 5'b01111; w[14][31] = 5'b00000; w[14][32] = 5'b10000; w[14][33] = 5'b10000; w[14][34] = 5'b10000; w[14][35] = 5'b10000; w[14][36] = 5'b10000; w[14][37] = 5'b10000; w[14][38] = 5'b00000; w[14][39] = 5'b01111; w[14][40] = 5'b01111; w[14][41] = 5'b01111; w[14][42] = 5'b01111; w[14][43] = 5'b01111; w[14][44] = 5'b01111; w[14][45] = 5'b10000; w[14][46] = 5'b10000; w[14][47] = 5'b10000; w[14][48] = 5'b10000; w[14][49] = 5'b10000; w[14][50] = 5'b10000; w[14][51] = 5'b10000; w[14][52] = 5'b10000; w[14][53] = 5'b01111; w[14][54] = 5'b01111; w[14][55] = 5'b01111; w[14][56] = 5'b01111; w[14][57] = 5'b01111; w[14][58] = 5'b01111; w[14][59] = 5'b00000; w[14][60] = 5'b00000; w[14][61] = 5'b01111; w[14][62] = 5'b10000; w[14][63] = 5'b00000; w[14][64] = 5'b01111; w[14][65] = 5'b00000; w[14][66] = 5'b00000; w[14][67] = 5'b01111; w[14][68] = 5'b01111; w[14][69] = 5'b01111; w[14][70] = 5'b01111; w[14][71] = 5'b01111; w[14][72] = 5'b01111; w[14][73] = 5'b00000; w[14][74] = 5'b01111; w[14][75] = 5'b01111; w[14][76] = 5'b10000; w[14][77] = 5'b00000; w[14][78] = 5'b01111; w[14][79] = 5'b01111; w[14][80] = 5'b00000; w[14][81] = 5'b01111; w[14][82] = 5'b01111; w[14][83] = 5'b01111; w[14][84] = 5'b01111; w[14][85] = 5'b01111; w[14][86] = 5'b01111; w[14][87] = 5'b00000; w[14][88] = 5'b01111; w[14][89] = 5'b01111; w[14][90] = 5'b10000; w[14][91] = 5'b10000; w[14][92] = 5'b01111; w[14][93] = 5'b01111; w[14][94] = 5'b01111; w[14][95] = 5'b01111; w[14][96] = 5'b01111; w[14][97] = 5'b01111; w[14][98] = 5'b01111; w[14][99] = 5'b01111; w[14][100] = 5'b01111; w[14][101] = 5'b00000; w[14][102] = 5'b01111; w[14][103] = 5'b01111; w[14][104] = 5'b10000; w[14][105] = 5'b10000; w[14][106] = 5'b01111; w[14][107] = 5'b00000; w[14][108] = 5'b00000; w[14][109] = 5'b01111; w[14][110] = 5'b01111; w[14][111] = 5'b01111; w[14][112] = 5'b01111; w[14][113] = 5'b01111; w[14][114] = 5'b01111; w[14][115] = 5'b00000; w[14][116] = 5'b01111; w[14][117] = 5'b01111; w[14][118] = 5'b10000; w[14][119] = 5'b10000; w[14][120] = 5'b00000; w[14][121] = 5'b00000; w[14][122] = 5'b00000; w[14][123] = 5'b01111; w[14][124] = 5'b01111; w[14][125] = 5'b01111; w[14][126] = 5'b01111; w[14][127] = 5'b01111; w[14][128] = 5'b01111; w[14][129] = 5'b00000; w[14][130] = 5'b01111; w[14][131] = 5'b01111; w[14][132] = 5'b00000; w[14][133] = 5'b10000; w[14][134] = 5'b01111; w[14][135] = 5'b01111; w[14][136] = 5'b00000; w[14][137] = 5'b01111; w[14][138] = 5'b01111; w[14][139] = 5'b01111; w[14][140] = 5'b01111; w[14][141] = 5'b01111; w[14][142] = 5'b01111; w[14][143] = 5'b00000; w[14][144] = 5'b00000; w[14][145] = 5'b01111; w[14][146] = 5'b00000; w[14][147] = 5'b10000; w[14][148] = 5'b01111; w[14][149] = 5'b00000; w[14][150] = 5'b00000; w[14][151] = 5'b01111; w[14][152] = 5'b01111; w[14][153] = 5'b01111; w[14][154] = 5'b01111; w[14][155] = 5'b01111; w[14][156] = 5'b01111; w[14][157] = 5'b00000; w[14][158] = 5'b00000; w[14][159] = 5'b00000; w[14][160] = 5'b10000; w[14][161] = 5'b10000; w[14][162] = 5'b10000; w[14][163] = 5'b00000; w[14][164] = 5'b00000; w[14][165] = 5'b01111; w[14][166] = 5'b01111; w[14][167] = 5'b01111; w[14][168] = 5'b01111; w[14][169] = 5'b01111; w[14][170] = 5'b01111; w[14][171] = 5'b01111; w[14][172] = 5'b00000; w[14][173] = 5'b00000; w[14][174] = 5'b10000; w[14][175] = 5'b10000; w[14][176] = 5'b10000; w[14][177] = 5'b00000; w[14][178] = 5'b01111; w[14][179] = 5'b01111; w[14][180] = 5'b01111; w[14][181] = 5'b01111; w[14][182] = 5'b01111; w[14][183] = 5'b01111; w[14][184] = 5'b01111; w[14][185] = 5'b01111; w[14][186] = 5'b01111; w[14][187] = 5'b01111; w[14][188] = 5'b01111; w[14][189] = 5'b01111; w[14][190] = 5'b01111; w[14][191] = 5'b01111; w[14][192] = 5'b01111; w[14][193] = 5'b01111; w[14][194] = 5'b01111; w[14][195] = 5'b01111; w[14][196] = 5'b01111; w[14][197] = 5'b01111; w[14][198] = 5'b01111; w[14][199] = 5'b01111; w[14][200] = 5'b01111; w[14][201] = 5'b01111; w[14][202] = 5'b01111; w[14][203] = 5'b01111; w[14][204] = 5'b01111; w[14][205] = 5'b01111; w[14][206] = 5'b01111; w[14][207] = 5'b01111; w[14][208] = 5'b01111; w[14][209] = 5'b01111; 
w[15][0] = 5'b01111; w[15][1] = 5'b01111; w[15][2] = 5'b01111; w[15][3] = 5'b01111; w[15][4] = 5'b01111; w[15][5] = 5'b01111; w[15][6] = 5'b01111; w[15][7] = 5'b01111; w[15][8] = 5'b01111; w[15][9] = 5'b01111; w[15][10] = 5'b01111; w[15][11] = 5'b01111; w[15][12] = 5'b01111; w[15][13] = 5'b01111; w[15][14] = 5'b01111; w[15][15] = 5'b00000; w[15][16] = 5'b01111; w[15][17] = 5'b01111; w[15][18] = 5'b01111; w[15][19] = 5'b01111; w[15][20] = 5'b01111; w[15][21] = 5'b01111; w[15][22] = 5'b01111; w[15][23] = 5'b01111; w[15][24] = 5'b01111; w[15][25] = 5'b01111; w[15][26] = 5'b01111; w[15][27] = 5'b01111; w[15][28] = 5'b01111; w[15][29] = 5'b01111; w[15][30] = 5'b01111; w[15][31] = 5'b00000; w[15][32] = 5'b10000; w[15][33] = 5'b10000; w[15][34] = 5'b10000; w[15][35] = 5'b10000; w[15][36] = 5'b10000; w[15][37] = 5'b10000; w[15][38] = 5'b00000; w[15][39] = 5'b01111; w[15][40] = 5'b01111; w[15][41] = 5'b01111; w[15][42] = 5'b01111; w[15][43] = 5'b01111; w[15][44] = 5'b01111; w[15][45] = 5'b10000; w[15][46] = 5'b10000; w[15][47] = 5'b10000; w[15][48] = 5'b10000; w[15][49] = 5'b10000; w[15][50] = 5'b10000; w[15][51] = 5'b10000; w[15][52] = 5'b10000; w[15][53] = 5'b01111; w[15][54] = 5'b01111; w[15][55] = 5'b01111; w[15][56] = 5'b01111; w[15][57] = 5'b01111; w[15][58] = 5'b01111; w[15][59] = 5'b00000; w[15][60] = 5'b00000; w[15][61] = 5'b01111; w[15][62] = 5'b10000; w[15][63] = 5'b00000; w[15][64] = 5'b01111; w[15][65] = 5'b00000; w[15][66] = 5'b00000; w[15][67] = 5'b01111; w[15][68] = 5'b01111; w[15][69] = 5'b01111; w[15][70] = 5'b01111; w[15][71] = 5'b01111; w[15][72] = 5'b01111; w[15][73] = 5'b00000; w[15][74] = 5'b01111; w[15][75] = 5'b01111; w[15][76] = 5'b10000; w[15][77] = 5'b00000; w[15][78] = 5'b01111; w[15][79] = 5'b01111; w[15][80] = 5'b00000; w[15][81] = 5'b01111; w[15][82] = 5'b01111; w[15][83] = 5'b01111; w[15][84] = 5'b01111; w[15][85] = 5'b01111; w[15][86] = 5'b01111; w[15][87] = 5'b00000; w[15][88] = 5'b01111; w[15][89] = 5'b01111; w[15][90] = 5'b10000; w[15][91] = 5'b10000; w[15][92] = 5'b01111; w[15][93] = 5'b01111; w[15][94] = 5'b01111; w[15][95] = 5'b01111; w[15][96] = 5'b01111; w[15][97] = 5'b01111; w[15][98] = 5'b01111; w[15][99] = 5'b01111; w[15][100] = 5'b01111; w[15][101] = 5'b00000; w[15][102] = 5'b01111; w[15][103] = 5'b01111; w[15][104] = 5'b10000; w[15][105] = 5'b10000; w[15][106] = 5'b01111; w[15][107] = 5'b00000; w[15][108] = 5'b00000; w[15][109] = 5'b01111; w[15][110] = 5'b01111; w[15][111] = 5'b01111; w[15][112] = 5'b01111; w[15][113] = 5'b01111; w[15][114] = 5'b01111; w[15][115] = 5'b00000; w[15][116] = 5'b01111; w[15][117] = 5'b01111; w[15][118] = 5'b10000; w[15][119] = 5'b10000; w[15][120] = 5'b00000; w[15][121] = 5'b00000; w[15][122] = 5'b00000; w[15][123] = 5'b01111; w[15][124] = 5'b01111; w[15][125] = 5'b01111; w[15][126] = 5'b01111; w[15][127] = 5'b01111; w[15][128] = 5'b01111; w[15][129] = 5'b00000; w[15][130] = 5'b01111; w[15][131] = 5'b01111; w[15][132] = 5'b00000; w[15][133] = 5'b10000; w[15][134] = 5'b01111; w[15][135] = 5'b01111; w[15][136] = 5'b00000; w[15][137] = 5'b01111; w[15][138] = 5'b01111; w[15][139] = 5'b01111; w[15][140] = 5'b01111; w[15][141] = 5'b01111; w[15][142] = 5'b01111; w[15][143] = 5'b00000; w[15][144] = 5'b00000; w[15][145] = 5'b01111; w[15][146] = 5'b00000; w[15][147] = 5'b10000; w[15][148] = 5'b01111; w[15][149] = 5'b00000; w[15][150] = 5'b00000; w[15][151] = 5'b01111; w[15][152] = 5'b01111; w[15][153] = 5'b01111; w[15][154] = 5'b01111; w[15][155] = 5'b01111; w[15][156] = 5'b01111; w[15][157] = 5'b00000; w[15][158] = 5'b00000; w[15][159] = 5'b00000; w[15][160] = 5'b10000; w[15][161] = 5'b10000; w[15][162] = 5'b10000; w[15][163] = 5'b00000; w[15][164] = 5'b00000; w[15][165] = 5'b01111; w[15][166] = 5'b01111; w[15][167] = 5'b01111; w[15][168] = 5'b01111; w[15][169] = 5'b01111; w[15][170] = 5'b01111; w[15][171] = 5'b01111; w[15][172] = 5'b00000; w[15][173] = 5'b00000; w[15][174] = 5'b10000; w[15][175] = 5'b10000; w[15][176] = 5'b10000; w[15][177] = 5'b00000; w[15][178] = 5'b01111; w[15][179] = 5'b01111; w[15][180] = 5'b01111; w[15][181] = 5'b01111; w[15][182] = 5'b01111; w[15][183] = 5'b01111; w[15][184] = 5'b01111; w[15][185] = 5'b01111; w[15][186] = 5'b01111; w[15][187] = 5'b01111; w[15][188] = 5'b01111; w[15][189] = 5'b01111; w[15][190] = 5'b01111; w[15][191] = 5'b01111; w[15][192] = 5'b01111; w[15][193] = 5'b01111; w[15][194] = 5'b01111; w[15][195] = 5'b01111; w[15][196] = 5'b01111; w[15][197] = 5'b01111; w[15][198] = 5'b01111; w[15][199] = 5'b01111; w[15][200] = 5'b01111; w[15][201] = 5'b01111; w[15][202] = 5'b01111; w[15][203] = 5'b01111; w[15][204] = 5'b01111; w[15][205] = 5'b01111; w[15][206] = 5'b01111; w[15][207] = 5'b01111; w[15][208] = 5'b01111; w[15][209] = 5'b01111; 
w[16][0] = 5'b01111; w[16][1] = 5'b01111; w[16][2] = 5'b01111; w[16][3] = 5'b01111; w[16][4] = 5'b01111; w[16][5] = 5'b01111; w[16][6] = 5'b01111; w[16][7] = 5'b01111; w[16][8] = 5'b01111; w[16][9] = 5'b01111; w[16][10] = 5'b01111; w[16][11] = 5'b01111; w[16][12] = 5'b01111; w[16][13] = 5'b01111; w[16][14] = 5'b01111; w[16][15] = 5'b01111; w[16][16] = 5'b00000; w[16][17] = 5'b01111; w[16][18] = 5'b01111; w[16][19] = 5'b01111; w[16][20] = 5'b01111; w[16][21] = 5'b01111; w[16][22] = 5'b01111; w[16][23] = 5'b01111; w[16][24] = 5'b01111; w[16][25] = 5'b01111; w[16][26] = 5'b01111; w[16][27] = 5'b01111; w[16][28] = 5'b01111; w[16][29] = 5'b01111; w[16][30] = 5'b01111; w[16][31] = 5'b00000; w[16][32] = 5'b10000; w[16][33] = 5'b10000; w[16][34] = 5'b10000; w[16][35] = 5'b10000; w[16][36] = 5'b10000; w[16][37] = 5'b10000; w[16][38] = 5'b00000; w[16][39] = 5'b01111; w[16][40] = 5'b01111; w[16][41] = 5'b01111; w[16][42] = 5'b01111; w[16][43] = 5'b01111; w[16][44] = 5'b01111; w[16][45] = 5'b10000; w[16][46] = 5'b10000; w[16][47] = 5'b10000; w[16][48] = 5'b10000; w[16][49] = 5'b10000; w[16][50] = 5'b10000; w[16][51] = 5'b10000; w[16][52] = 5'b10000; w[16][53] = 5'b01111; w[16][54] = 5'b01111; w[16][55] = 5'b01111; w[16][56] = 5'b01111; w[16][57] = 5'b01111; w[16][58] = 5'b01111; w[16][59] = 5'b00000; w[16][60] = 5'b00000; w[16][61] = 5'b01111; w[16][62] = 5'b10000; w[16][63] = 5'b00000; w[16][64] = 5'b01111; w[16][65] = 5'b00000; w[16][66] = 5'b00000; w[16][67] = 5'b01111; w[16][68] = 5'b01111; w[16][69] = 5'b01111; w[16][70] = 5'b01111; w[16][71] = 5'b01111; w[16][72] = 5'b01111; w[16][73] = 5'b00000; w[16][74] = 5'b01111; w[16][75] = 5'b01111; w[16][76] = 5'b10000; w[16][77] = 5'b00000; w[16][78] = 5'b01111; w[16][79] = 5'b01111; w[16][80] = 5'b00000; w[16][81] = 5'b01111; w[16][82] = 5'b01111; w[16][83] = 5'b01111; w[16][84] = 5'b01111; w[16][85] = 5'b01111; w[16][86] = 5'b01111; w[16][87] = 5'b00000; w[16][88] = 5'b01111; w[16][89] = 5'b01111; w[16][90] = 5'b10000; w[16][91] = 5'b10000; w[16][92] = 5'b01111; w[16][93] = 5'b01111; w[16][94] = 5'b01111; w[16][95] = 5'b01111; w[16][96] = 5'b01111; w[16][97] = 5'b01111; w[16][98] = 5'b01111; w[16][99] = 5'b01111; w[16][100] = 5'b01111; w[16][101] = 5'b00000; w[16][102] = 5'b01111; w[16][103] = 5'b01111; w[16][104] = 5'b10000; w[16][105] = 5'b10000; w[16][106] = 5'b01111; w[16][107] = 5'b00000; w[16][108] = 5'b00000; w[16][109] = 5'b01111; w[16][110] = 5'b01111; w[16][111] = 5'b01111; w[16][112] = 5'b01111; w[16][113] = 5'b01111; w[16][114] = 5'b01111; w[16][115] = 5'b00000; w[16][116] = 5'b01111; w[16][117] = 5'b01111; w[16][118] = 5'b10000; w[16][119] = 5'b10000; w[16][120] = 5'b00000; w[16][121] = 5'b00000; w[16][122] = 5'b00000; w[16][123] = 5'b01111; w[16][124] = 5'b01111; w[16][125] = 5'b01111; w[16][126] = 5'b01111; w[16][127] = 5'b01111; w[16][128] = 5'b01111; w[16][129] = 5'b00000; w[16][130] = 5'b01111; w[16][131] = 5'b01111; w[16][132] = 5'b00000; w[16][133] = 5'b10000; w[16][134] = 5'b01111; w[16][135] = 5'b01111; w[16][136] = 5'b00000; w[16][137] = 5'b01111; w[16][138] = 5'b01111; w[16][139] = 5'b01111; w[16][140] = 5'b01111; w[16][141] = 5'b01111; w[16][142] = 5'b01111; w[16][143] = 5'b00000; w[16][144] = 5'b00000; w[16][145] = 5'b01111; w[16][146] = 5'b00000; w[16][147] = 5'b10000; w[16][148] = 5'b01111; w[16][149] = 5'b00000; w[16][150] = 5'b00000; w[16][151] = 5'b01111; w[16][152] = 5'b01111; w[16][153] = 5'b01111; w[16][154] = 5'b01111; w[16][155] = 5'b01111; w[16][156] = 5'b01111; w[16][157] = 5'b00000; w[16][158] = 5'b00000; w[16][159] = 5'b00000; w[16][160] = 5'b10000; w[16][161] = 5'b10000; w[16][162] = 5'b10000; w[16][163] = 5'b00000; w[16][164] = 5'b00000; w[16][165] = 5'b01111; w[16][166] = 5'b01111; w[16][167] = 5'b01111; w[16][168] = 5'b01111; w[16][169] = 5'b01111; w[16][170] = 5'b01111; w[16][171] = 5'b01111; w[16][172] = 5'b00000; w[16][173] = 5'b00000; w[16][174] = 5'b10000; w[16][175] = 5'b10000; w[16][176] = 5'b10000; w[16][177] = 5'b00000; w[16][178] = 5'b01111; w[16][179] = 5'b01111; w[16][180] = 5'b01111; w[16][181] = 5'b01111; w[16][182] = 5'b01111; w[16][183] = 5'b01111; w[16][184] = 5'b01111; w[16][185] = 5'b01111; w[16][186] = 5'b01111; w[16][187] = 5'b01111; w[16][188] = 5'b01111; w[16][189] = 5'b01111; w[16][190] = 5'b01111; w[16][191] = 5'b01111; w[16][192] = 5'b01111; w[16][193] = 5'b01111; w[16][194] = 5'b01111; w[16][195] = 5'b01111; w[16][196] = 5'b01111; w[16][197] = 5'b01111; w[16][198] = 5'b01111; w[16][199] = 5'b01111; w[16][200] = 5'b01111; w[16][201] = 5'b01111; w[16][202] = 5'b01111; w[16][203] = 5'b01111; w[16][204] = 5'b01111; w[16][205] = 5'b01111; w[16][206] = 5'b01111; w[16][207] = 5'b01111; w[16][208] = 5'b01111; w[16][209] = 5'b01111; 
w[17][0] = 5'b01111; w[17][1] = 5'b01111; w[17][2] = 5'b01111; w[17][3] = 5'b01111; w[17][4] = 5'b01111; w[17][5] = 5'b01111; w[17][6] = 5'b01111; w[17][7] = 5'b01111; w[17][8] = 5'b01111; w[17][9] = 5'b01111; w[17][10] = 5'b01111; w[17][11] = 5'b01111; w[17][12] = 5'b01111; w[17][13] = 5'b01111; w[17][14] = 5'b01111; w[17][15] = 5'b01111; w[17][16] = 5'b01111; w[17][17] = 5'b00000; w[17][18] = 5'b01111; w[17][19] = 5'b01111; w[17][20] = 5'b01111; w[17][21] = 5'b01111; w[17][22] = 5'b01111; w[17][23] = 5'b01111; w[17][24] = 5'b01111; w[17][25] = 5'b01111; w[17][26] = 5'b01111; w[17][27] = 5'b01111; w[17][28] = 5'b01111; w[17][29] = 5'b01111; w[17][30] = 5'b01111; w[17][31] = 5'b00000; w[17][32] = 5'b10000; w[17][33] = 5'b10000; w[17][34] = 5'b10000; w[17][35] = 5'b10000; w[17][36] = 5'b10000; w[17][37] = 5'b10000; w[17][38] = 5'b00000; w[17][39] = 5'b01111; w[17][40] = 5'b01111; w[17][41] = 5'b01111; w[17][42] = 5'b01111; w[17][43] = 5'b01111; w[17][44] = 5'b01111; w[17][45] = 5'b10000; w[17][46] = 5'b10000; w[17][47] = 5'b10000; w[17][48] = 5'b10000; w[17][49] = 5'b10000; w[17][50] = 5'b10000; w[17][51] = 5'b10000; w[17][52] = 5'b10000; w[17][53] = 5'b01111; w[17][54] = 5'b01111; w[17][55] = 5'b01111; w[17][56] = 5'b01111; w[17][57] = 5'b01111; w[17][58] = 5'b01111; w[17][59] = 5'b00000; w[17][60] = 5'b00000; w[17][61] = 5'b01111; w[17][62] = 5'b10000; w[17][63] = 5'b00000; w[17][64] = 5'b01111; w[17][65] = 5'b00000; w[17][66] = 5'b00000; w[17][67] = 5'b01111; w[17][68] = 5'b01111; w[17][69] = 5'b01111; w[17][70] = 5'b01111; w[17][71] = 5'b01111; w[17][72] = 5'b01111; w[17][73] = 5'b00000; w[17][74] = 5'b01111; w[17][75] = 5'b01111; w[17][76] = 5'b10000; w[17][77] = 5'b00000; w[17][78] = 5'b01111; w[17][79] = 5'b01111; w[17][80] = 5'b00000; w[17][81] = 5'b01111; w[17][82] = 5'b01111; w[17][83] = 5'b01111; w[17][84] = 5'b01111; w[17][85] = 5'b01111; w[17][86] = 5'b01111; w[17][87] = 5'b00000; w[17][88] = 5'b01111; w[17][89] = 5'b01111; w[17][90] = 5'b10000; w[17][91] = 5'b10000; w[17][92] = 5'b01111; w[17][93] = 5'b01111; w[17][94] = 5'b01111; w[17][95] = 5'b01111; w[17][96] = 5'b01111; w[17][97] = 5'b01111; w[17][98] = 5'b01111; w[17][99] = 5'b01111; w[17][100] = 5'b01111; w[17][101] = 5'b00000; w[17][102] = 5'b01111; w[17][103] = 5'b01111; w[17][104] = 5'b10000; w[17][105] = 5'b10000; w[17][106] = 5'b01111; w[17][107] = 5'b00000; w[17][108] = 5'b00000; w[17][109] = 5'b01111; w[17][110] = 5'b01111; w[17][111] = 5'b01111; w[17][112] = 5'b01111; w[17][113] = 5'b01111; w[17][114] = 5'b01111; w[17][115] = 5'b00000; w[17][116] = 5'b01111; w[17][117] = 5'b01111; w[17][118] = 5'b10000; w[17][119] = 5'b10000; w[17][120] = 5'b00000; w[17][121] = 5'b00000; w[17][122] = 5'b00000; w[17][123] = 5'b01111; w[17][124] = 5'b01111; w[17][125] = 5'b01111; w[17][126] = 5'b01111; w[17][127] = 5'b01111; w[17][128] = 5'b01111; w[17][129] = 5'b00000; w[17][130] = 5'b01111; w[17][131] = 5'b01111; w[17][132] = 5'b00000; w[17][133] = 5'b10000; w[17][134] = 5'b01111; w[17][135] = 5'b01111; w[17][136] = 5'b00000; w[17][137] = 5'b01111; w[17][138] = 5'b01111; w[17][139] = 5'b01111; w[17][140] = 5'b01111; w[17][141] = 5'b01111; w[17][142] = 5'b01111; w[17][143] = 5'b00000; w[17][144] = 5'b00000; w[17][145] = 5'b01111; w[17][146] = 5'b00000; w[17][147] = 5'b10000; w[17][148] = 5'b01111; w[17][149] = 5'b00000; w[17][150] = 5'b00000; w[17][151] = 5'b01111; w[17][152] = 5'b01111; w[17][153] = 5'b01111; w[17][154] = 5'b01111; w[17][155] = 5'b01111; w[17][156] = 5'b01111; w[17][157] = 5'b00000; w[17][158] = 5'b00000; w[17][159] = 5'b00000; w[17][160] = 5'b10000; w[17][161] = 5'b10000; w[17][162] = 5'b10000; w[17][163] = 5'b00000; w[17][164] = 5'b00000; w[17][165] = 5'b01111; w[17][166] = 5'b01111; w[17][167] = 5'b01111; w[17][168] = 5'b01111; w[17][169] = 5'b01111; w[17][170] = 5'b01111; w[17][171] = 5'b01111; w[17][172] = 5'b00000; w[17][173] = 5'b00000; w[17][174] = 5'b10000; w[17][175] = 5'b10000; w[17][176] = 5'b10000; w[17][177] = 5'b00000; w[17][178] = 5'b01111; w[17][179] = 5'b01111; w[17][180] = 5'b01111; w[17][181] = 5'b01111; w[17][182] = 5'b01111; w[17][183] = 5'b01111; w[17][184] = 5'b01111; w[17][185] = 5'b01111; w[17][186] = 5'b01111; w[17][187] = 5'b01111; w[17][188] = 5'b01111; w[17][189] = 5'b01111; w[17][190] = 5'b01111; w[17][191] = 5'b01111; w[17][192] = 5'b01111; w[17][193] = 5'b01111; w[17][194] = 5'b01111; w[17][195] = 5'b01111; w[17][196] = 5'b01111; w[17][197] = 5'b01111; w[17][198] = 5'b01111; w[17][199] = 5'b01111; w[17][200] = 5'b01111; w[17][201] = 5'b01111; w[17][202] = 5'b01111; w[17][203] = 5'b01111; w[17][204] = 5'b01111; w[17][205] = 5'b01111; w[17][206] = 5'b01111; w[17][207] = 5'b01111; w[17][208] = 5'b01111; w[17][209] = 5'b01111; 
w[18][0] = 5'b01111; w[18][1] = 5'b01111; w[18][2] = 5'b01111; w[18][3] = 5'b01111; w[18][4] = 5'b01111; w[18][5] = 5'b01111; w[18][6] = 5'b01111; w[18][7] = 5'b01111; w[18][8] = 5'b01111; w[18][9] = 5'b01111; w[18][10] = 5'b01111; w[18][11] = 5'b01111; w[18][12] = 5'b01111; w[18][13] = 5'b01111; w[18][14] = 5'b01111; w[18][15] = 5'b01111; w[18][16] = 5'b01111; w[18][17] = 5'b01111; w[18][18] = 5'b00000; w[18][19] = 5'b01111; w[18][20] = 5'b01111; w[18][21] = 5'b01111; w[18][22] = 5'b01111; w[18][23] = 5'b01111; w[18][24] = 5'b01111; w[18][25] = 5'b01111; w[18][26] = 5'b01111; w[18][27] = 5'b01111; w[18][28] = 5'b01111; w[18][29] = 5'b01111; w[18][30] = 5'b01111; w[18][31] = 5'b00000; w[18][32] = 5'b10000; w[18][33] = 5'b10000; w[18][34] = 5'b10000; w[18][35] = 5'b10000; w[18][36] = 5'b10000; w[18][37] = 5'b10000; w[18][38] = 5'b00000; w[18][39] = 5'b01111; w[18][40] = 5'b01111; w[18][41] = 5'b01111; w[18][42] = 5'b01111; w[18][43] = 5'b01111; w[18][44] = 5'b01111; w[18][45] = 5'b10000; w[18][46] = 5'b10000; w[18][47] = 5'b10000; w[18][48] = 5'b10000; w[18][49] = 5'b10000; w[18][50] = 5'b10000; w[18][51] = 5'b10000; w[18][52] = 5'b10000; w[18][53] = 5'b01111; w[18][54] = 5'b01111; w[18][55] = 5'b01111; w[18][56] = 5'b01111; w[18][57] = 5'b01111; w[18][58] = 5'b01111; w[18][59] = 5'b00000; w[18][60] = 5'b00000; w[18][61] = 5'b01111; w[18][62] = 5'b10000; w[18][63] = 5'b00000; w[18][64] = 5'b01111; w[18][65] = 5'b00000; w[18][66] = 5'b00000; w[18][67] = 5'b01111; w[18][68] = 5'b01111; w[18][69] = 5'b01111; w[18][70] = 5'b01111; w[18][71] = 5'b01111; w[18][72] = 5'b01111; w[18][73] = 5'b00000; w[18][74] = 5'b01111; w[18][75] = 5'b01111; w[18][76] = 5'b10000; w[18][77] = 5'b00000; w[18][78] = 5'b01111; w[18][79] = 5'b01111; w[18][80] = 5'b00000; w[18][81] = 5'b01111; w[18][82] = 5'b01111; w[18][83] = 5'b01111; w[18][84] = 5'b01111; w[18][85] = 5'b01111; w[18][86] = 5'b01111; w[18][87] = 5'b00000; w[18][88] = 5'b01111; w[18][89] = 5'b01111; w[18][90] = 5'b10000; w[18][91] = 5'b10000; w[18][92] = 5'b01111; w[18][93] = 5'b01111; w[18][94] = 5'b01111; w[18][95] = 5'b01111; w[18][96] = 5'b01111; w[18][97] = 5'b01111; w[18][98] = 5'b01111; w[18][99] = 5'b01111; w[18][100] = 5'b01111; w[18][101] = 5'b00000; w[18][102] = 5'b01111; w[18][103] = 5'b01111; w[18][104] = 5'b10000; w[18][105] = 5'b10000; w[18][106] = 5'b01111; w[18][107] = 5'b00000; w[18][108] = 5'b00000; w[18][109] = 5'b01111; w[18][110] = 5'b01111; w[18][111] = 5'b01111; w[18][112] = 5'b01111; w[18][113] = 5'b01111; w[18][114] = 5'b01111; w[18][115] = 5'b00000; w[18][116] = 5'b01111; w[18][117] = 5'b01111; w[18][118] = 5'b10000; w[18][119] = 5'b10000; w[18][120] = 5'b00000; w[18][121] = 5'b00000; w[18][122] = 5'b00000; w[18][123] = 5'b01111; w[18][124] = 5'b01111; w[18][125] = 5'b01111; w[18][126] = 5'b01111; w[18][127] = 5'b01111; w[18][128] = 5'b01111; w[18][129] = 5'b00000; w[18][130] = 5'b01111; w[18][131] = 5'b01111; w[18][132] = 5'b00000; w[18][133] = 5'b10000; w[18][134] = 5'b01111; w[18][135] = 5'b01111; w[18][136] = 5'b00000; w[18][137] = 5'b01111; w[18][138] = 5'b01111; w[18][139] = 5'b01111; w[18][140] = 5'b01111; w[18][141] = 5'b01111; w[18][142] = 5'b01111; w[18][143] = 5'b00000; w[18][144] = 5'b00000; w[18][145] = 5'b01111; w[18][146] = 5'b00000; w[18][147] = 5'b10000; w[18][148] = 5'b01111; w[18][149] = 5'b00000; w[18][150] = 5'b00000; w[18][151] = 5'b01111; w[18][152] = 5'b01111; w[18][153] = 5'b01111; w[18][154] = 5'b01111; w[18][155] = 5'b01111; w[18][156] = 5'b01111; w[18][157] = 5'b00000; w[18][158] = 5'b00000; w[18][159] = 5'b00000; w[18][160] = 5'b10000; w[18][161] = 5'b10000; w[18][162] = 5'b10000; w[18][163] = 5'b00000; w[18][164] = 5'b00000; w[18][165] = 5'b01111; w[18][166] = 5'b01111; w[18][167] = 5'b01111; w[18][168] = 5'b01111; w[18][169] = 5'b01111; w[18][170] = 5'b01111; w[18][171] = 5'b01111; w[18][172] = 5'b00000; w[18][173] = 5'b00000; w[18][174] = 5'b10000; w[18][175] = 5'b10000; w[18][176] = 5'b10000; w[18][177] = 5'b00000; w[18][178] = 5'b01111; w[18][179] = 5'b01111; w[18][180] = 5'b01111; w[18][181] = 5'b01111; w[18][182] = 5'b01111; w[18][183] = 5'b01111; w[18][184] = 5'b01111; w[18][185] = 5'b01111; w[18][186] = 5'b01111; w[18][187] = 5'b01111; w[18][188] = 5'b01111; w[18][189] = 5'b01111; w[18][190] = 5'b01111; w[18][191] = 5'b01111; w[18][192] = 5'b01111; w[18][193] = 5'b01111; w[18][194] = 5'b01111; w[18][195] = 5'b01111; w[18][196] = 5'b01111; w[18][197] = 5'b01111; w[18][198] = 5'b01111; w[18][199] = 5'b01111; w[18][200] = 5'b01111; w[18][201] = 5'b01111; w[18][202] = 5'b01111; w[18][203] = 5'b01111; w[18][204] = 5'b01111; w[18][205] = 5'b01111; w[18][206] = 5'b01111; w[18][207] = 5'b01111; w[18][208] = 5'b01111; w[18][209] = 5'b01111; 
w[19][0] = 5'b01111; w[19][1] = 5'b01111; w[19][2] = 5'b01111; w[19][3] = 5'b01111; w[19][4] = 5'b01111; w[19][5] = 5'b01111; w[19][6] = 5'b01111; w[19][7] = 5'b01111; w[19][8] = 5'b01111; w[19][9] = 5'b01111; w[19][10] = 5'b01111; w[19][11] = 5'b01111; w[19][12] = 5'b01111; w[19][13] = 5'b01111; w[19][14] = 5'b01111; w[19][15] = 5'b01111; w[19][16] = 5'b01111; w[19][17] = 5'b01111; w[19][18] = 5'b01111; w[19][19] = 5'b00000; w[19][20] = 5'b01111; w[19][21] = 5'b01111; w[19][22] = 5'b01111; w[19][23] = 5'b01111; w[19][24] = 5'b01111; w[19][25] = 5'b01111; w[19][26] = 5'b01111; w[19][27] = 5'b01111; w[19][28] = 5'b01111; w[19][29] = 5'b01111; w[19][30] = 5'b01111; w[19][31] = 5'b00000; w[19][32] = 5'b10000; w[19][33] = 5'b10000; w[19][34] = 5'b10000; w[19][35] = 5'b10000; w[19][36] = 5'b10000; w[19][37] = 5'b10000; w[19][38] = 5'b00000; w[19][39] = 5'b01111; w[19][40] = 5'b01111; w[19][41] = 5'b01111; w[19][42] = 5'b01111; w[19][43] = 5'b01111; w[19][44] = 5'b01111; w[19][45] = 5'b10000; w[19][46] = 5'b10000; w[19][47] = 5'b10000; w[19][48] = 5'b10000; w[19][49] = 5'b10000; w[19][50] = 5'b10000; w[19][51] = 5'b10000; w[19][52] = 5'b10000; w[19][53] = 5'b01111; w[19][54] = 5'b01111; w[19][55] = 5'b01111; w[19][56] = 5'b01111; w[19][57] = 5'b01111; w[19][58] = 5'b01111; w[19][59] = 5'b00000; w[19][60] = 5'b00000; w[19][61] = 5'b01111; w[19][62] = 5'b10000; w[19][63] = 5'b00000; w[19][64] = 5'b01111; w[19][65] = 5'b00000; w[19][66] = 5'b00000; w[19][67] = 5'b01111; w[19][68] = 5'b01111; w[19][69] = 5'b01111; w[19][70] = 5'b01111; w[19][71] = 5'b01111; w[19][72] = 5'b01111; w[19][73] = 5'b00000; w[19][74] = 5'b01111; w[19][75] = 5'b01111; w[19][76] = 5'b10000; w[19][77] = 5'b00000; w[19][78] = 5'b01111; w[19][79] = 5'b01111; w[19][80] = 5'b00000; w[19][81] = 5'b01111; w[19][82] = 5'b01111; w[19][83] = 5'b01111; w[19][84] = 5'b01111; w[19][85] = 5'b01111; w[19][86] = 5'b01111; w[19][87] = 5'b00000; w[19][88] = 5'b01111; w[19][89] = 5'b01111; w[19][90] = 5'b10000; w[19][91] = 5'b10000; w[19][92] = 5'b01111; w[19][93] = 5'b01111; w[19][94] = 5'b01111; w[19][95] = 5'b01111; w[19][96] = 5'b01111; w[19][97] = 5'b01111; w[19][98] = 5'b01111; w[19][99] = 5'b01111; w[19][100] = 5'b01111; w[19][101] = 5'b00000; w[19][102] = 5'b01111; w[19][103] = 5'b01111; w[19][104] = 5'b10000; w[19][105] = 5'b10000; w[19][106] = 5'b01111; w[19][107] = 5'b00000; w[19][108] = 5'b00000; w[19][109] = 5'b01111; w[19][110] = 5'b01111; w[19][111] = 5'b01111; w[19][112] = 5'b01111; w[19][113] = 5'b01111; w[19][114] = 5'b01111; w[19][115] = 5'b00000; w[19][116] = 5'b01111; w[19][117] = 5'b01111; w[19][118] = 5'b10000; w[19][119] = 5'b10000; w[19][120] = 5'b00000; w[19][121] = 5'b00000; w[19][122] = 5'b00000; w[19][123] = 5'b01111; w[19][124] = 5'b01111; w[19][125] = 5'b01111; w[19][126] = 5'b01111; w[19][127] = 5'b01111; w[19][128] = 5'b01111; w[19][129] = 5'b00000; w[19][130] = 5'b01111; w[19][131] = 5'b01111; w[19][132] = 5'b00000; w[19][133] = 5'b10000; w[19][134] = 5'b01111; w[19][135] = 5'b01111; w[19][136] = 5'b00000; w[19][137] = 5'b01111; w[19][138] = 5'b01111; w[19][139] = 5'b01111; w[19][140] = 5'b01111; w[19][141] = 5'b01111; w[19][142] = 5'b01111; w[19][143] = 5'b00000; w[19][144] = 5'b00000; w[19][145] = 5'b01111; w[19][146] = 5'b00000; w[19][147] = 5'b10000; w[19][148] = 5'b01111; w[19][149] = 5'b00000; w[19][150] = 5'b00000; w[19][151] = 5'b01111; w[19][152] = 5'b01111; w[19][153] = 5'b01111; w[19][154] = 5'b01111; w[19][155] = 5'b01111; w[19][156] = 5'b01111; w[19][157] = 5'b00000; w[19][158] = 5'b00000; w[19][159] = 5'b00000; w[19][160] = 5'b10000; w[19][161] = 5'b10000; w[19][162] = 5'b10000; w[19][163] = 5'b00000; w[19][164] = 5'b00000; w[19][165] = 5'b01111; w[19][166] = 5'b01111; w[19][167] = 5'b01111; w[19][168] = 5'b01111; w[19][169] = 5'b01111; w[19][170] = 5'b01111; w[19][171] = 5'b01111; w[19][172] = 5'b00000; w[19][173] = 5'b00000; w[19][174] = 5'b10000; w[19][175] = 5'b10000; w[19][176] = 5'b10000; w[19][177] = 5'b00000; w[19][178] = 5'b01111; w[19][179] = 5'b01111; w[19][180] = 5'b01111; w[19][181] = 5'b01111; w[19][182] = 5'b01111; w[19][183] = 5'b01111; w[19][184] = 5'b01111; w[19][185] = 5'b01111; w[19][186] = 5'b01111; w[19][187] = 5'b01111; w[19][188] = 5'b01111; w[19][189] = 5'b01111; w[19][190] = 5'b01111; w[19][191] = 5'b01111; w[19][192] = 5'b01111; w[19][193] = 5'b01111; w[19][194] = 5'b01111; w[19][195] = 5'b01111; w[19][196] = 5'b01111; w[19][197] = 5'b01111; w[19][198] = 5'b01111; w[19][199] = 5'b01111; w[19][200] = 5'b01111; w[19][201] = 5'b01111; w[19][202] = 5'b01111; w[19][203] = 5'b01111; w[19][204] = 5'b01111; w[19][205] = 5'b01111; w[19][206] = 5'b01111; w[19][207] = 5'b01111; w[19][208] = 5'b01111; w[19][209] = 5'b01111; 
w[20][0] = 5'b01111; w[20][1] = 5'b01111; w[20][2] = 5'b01111; w[20][3] = 5'b01111; w[20][4] = 5'b01111; w[20][5] = 5'b01111; w[20][6] = 5'b01111; w[20][7] = 5'b01111; w[20][8] = 5'b01111; w[20][9] = 5'b01111; w[20][10] = 5'b01111; w[20][11] = 5'b01111; w[20][12] = 5'b01111; w[20][13] = 5'b01111; w[20][14] = 5'b01111; w[20][15] = 5'b01111; w[20][16] = 5'b01111; w[20][17] = 5'b01111; w[20][18] = 5'b01111; w[20][19] = 5'b01111; w[20][20] = 5'b00000; w[20][21] = 5'b01111; w[20][22] = 5'b01111; w[20][23] = 5'b01111; w[20][24] = 5'b01111; w[20][25] = 5'b01111; w[20][26] = 5'b01111; w[20][27] = 5'b01111; w[20][28] = 5'b01111; w[20][29] = 5'b01111; w[20][30] = 5'b01111; w[20][31] = 5'b00000; w[20][32] = 5'b10000; w[20][33] = 5'b10000; w[20][34] = 5'b10000; w[20][35] = 5'b10000; w[20][36] = 5'b10000; w[20][37] = 5'b10000; w[20][38] = 5'b00000; w[20][39] = 5'b01111; w[20][40] = 5'b01111; w[20][41] = 5'b01111; w[20][42] = 5'b01111; w[20][43] = 5'b01111; w[20][44] = 5'b01111; w[20][45] = 5'b10000; w[20][46] = 5'b10000; w[20][47] = 5'b10000; w[20][48] = 5'b10000; w[20][49] = 5'b10000; w[20][50] = 5'b10000; w[20][51] = 5'b10000; w[20][52] = 5'b10000; w[20][53] = 5'b01111; w[20][54] = 5'b01111; w[20][55] = 5'b01111; w[20][56] = 5'b01111; w[20][57] = 5'b01111; w[20][58] = 5'b01111; w[20][59] = 5'b00000; w[20][60] = 5'b00000; w[20][61] = 5'b01111; w[20][62] = 5'b10000; w[20][63] = 5'b00000; w[20][64] = 5'b01111; w[20][65] = 5'b00000; w[20][66] = 5'b00000; w[20][67] = 5'b01111; w[20][68] = 5'b01111; w[20][69] = 5'b01111; w[20][70] = 5'b01111; w[20][71] = 5'b01111; w[20][72] = 5'b01111; w[20][73] = 5'b00000; w[20][74] = 5'b01111; w[20][75] = 5'b01111; w[20][76] = 5'b10000; w[20][77] = 5'b00000; w[20][78] = 5'b01111; w[20][79] = 5'b01111; w[20][80] = 5'b00000; w[20][81] = 5'b01111; w[20][82] = 5'b01111; w[20][83] = 5'b01111; w[20][84] = 5'b01111; w[20][85] = 5'b01111; w[20][86] = 5'b01111; w[20][87] = 5'b00000; w[20][88] = 5'b01111; w[20][89] = 5'b01111; w[20][90] = 5'b10000; w[20][91] = 5'b10000; w[20][92] = 5'b01111; w[20][93] = 5'b01111; w[20][94] = 5'b01111; w[20][95] = 5'b01111; w[20][96] = 5'b01111; w[20][97] = 5'b01111; w[20][98] = 5'b01111; w[20][99] = 5'b01111; w[20][100] = 5'b01111; w[20][101] = 5'b00000; w[20][102] = 5'b01111; w[20][103] = 5'b01111; w[20][104] = 5'b10000; w[20][105] = 5'b10000; w[20][106] = 5'b01111; w[20][107] = 5'b00000; w[20][108] = 5'b00000; w[20][109] = 5'b01111; w[20][110] = 5'b01111; w[20][111] = 5'b01111; w[20][112] = 5'b01111; w[20][113] = 5'b01111; w[20][114] = 5'b01111; w[20][115] = 5'b00000; w[20][116] = 5'b01111; w[20][117] = 5'b01111; w[20][118] = 5'b10000; w[20][119] = 5'b10000; w[20][120] = 5'b00000; w[20][121] = 5'b00000; w[20][122] = 5'b00000; w[20][123] = 5'b01111; w[20][124] = 5'b01111; w[20][125] = 5'b01111; w[20][126] = 5'b01111; w[20][127] = 5'b01111; w[20][128] = 5'b01111; w[20][129] = 5'b00000; w[20][130] = 5'b01111; w[20][131] = 5'b01111; w[20][132] = 5'b00000; w[20][133] = 5'b10000; w[20][134] = 5'b01111; w[20][135] = 5'b01111; w[20][136] = 5'b00000; w[20][137] = 5'b01111; w[20][138] = 5'b01111; w[20][139] = 5'b01111; w[20][140] = 5'b01111; w[20][141] = 5'b01111; w[20][142] = 5'b01111; w[20][143] = 5'b00000; w[20][144] = 5'b00000; w[20][145] = 5'b01111; w[20][146] = 5'b00000; w[20][147] = 5'b10000; w[20][148] = 5'b01111; w[20][149] = 5'b00000; w[20][150] = 5'b00000; w[20][151] = 5'b01111; w[20][152] = 5'b01111; w[20][153] = 5'b01111; w[20][154] = 5'b01111; w[20][155] = 5'b01111; w[20][156] = 5'b01111; w[20][157] = 5'b00000; w[20][158] = 5'b00000; w[20][159] = 5'b00000; w[20][160] = 5'b10000; w[20][161] = 5'b10000; w[20][162] = 5'b10000; w[20][163] = 5'b00000; w[20][164] = 5'b00000; w[20][165] = 5'b01111; w[20][166] = 5'b01111; w[20][167] = 5'b01111; w[20][168] = 5'b01111; w[20][169] = 5'b01111; w[20][170] = 5'b01111; w[20][171] = 5'b01111; w[20][172] = 5'b00000; w[20][173] = 5'b00000; w[20][174] = 5'b10000; w[20][175] = 5'b10000; w[20][176] = 5'b10000; w[20][177] = 5'b00000; w[20][178] = 5'b01111; w[20][179] = 5'b01111; w[20][180] = 5'b01111; w[20][181] = 5'b01111; w[20][182] = 5'b01111; w[20][183] = 5'b01111; w[20][184] = 5'b01111; w[20][185] = 5'b01111; w[20][186] = 5'b01111; w[20][187] = 5'b01111; w[20][188] = 5'b01111; w[20][189] = 5'b01111; w[20][190] = 5'b01111; w[20][191] = 5'b01111; w[20][192] = 5'b01111; w[20][193] = 5'b01111; w[20][194] = 5'b01111; w[20][195] = 5'b01111; w[20][196] = 5'b01111; w[20][197] = 5'b01111; w[20][198] = 5'b01111; w[20][199] = 5'b01111; w[20][200] = 5'b01111; w[20][201] = 5'b01111; w[20][202] = 5'b01111; w[20][203] = 5'b01111; w[20][204] = 5'b01111; w[20][205] = 5'b01111; w[20][206] = 5'b01111; w[20][207] = 5'b01111; w[20][208] = 5'b01111; w[20][209] = 5'b01111; 
w[21][0] = 5'b01111; w[21][1] = 5'b01111; w[21][2] = 5'b01111; w[21][3] = 5'b01111; w[21][4] = 5'b01111; w[21][5] = 5'b01111; w[21][6] = 5'b01111; w[21][7] = 5'b01111; w[21][8] = 5'b01111; w[21][9] = 5'b01111; w[21][10] = 5'b01111; w[21][11] = 5'b01111; w[21][12] = 5'b01111; w[21][13] = 5'b01111; w[21][14] = 5'b01111; w[21][15] = 5'b01111; w[21][16] = 5'b01111; w[21][17] = 5'b01111; w[21][18] = 5'b01111; w[21][19] = 5'b01111; w[21][20] = 5'b01111; w[21][21] = 5'b00000; w[21][22] = 5'b01111; w[21][23] = 5'b01111; w[21][24] = 5'b01111; w[21][25] = 5'b01111; w[21][26] = 5'b01111; w[21][27] = 5'b01111; w[21][28] = 5'b01111; w[21][29] = 5'b01111; w[21][30] = 5'b01111; w[21][31] = 5'b00000; w[21][32] = 5'b10000; w[21][33] = 5'b10000; w[21][34] = 5'b10000; w[21][35] = 5'b10000; w[21][36] = 5'b10000; w[21][37] = 5'b10000; w[21][38] = 5'b00000; w[21][39] = 5'b01111; w[21][40] = 5'b01111; w[21][41] = 5'b01111; w[21][42] = 5'b01111; w[21][43] = 5'b01111; w[21][44] = 5'b01111; w[21][45] = 5'b10000; w[21][46] = 5'b10000; w[21][47] = 5'b10000; w[21][48] = 5'b10000; w[21][49] = 5'b10000; w[21][50] = 5'b10000; w[21][51] = 5'b10000; w[21][52] = 5'b10000; w[21][53] = 5'b01111; w[21][54] = 5'b01111; w[21][55] = 5'b01111; w[21][56] = 5'b01111; w[21][57] = 5'b01111; w[21][58] = 5'b01111; w[21][59] = 5'b00000; w[21][60] = 5'b00000; w[21][61] = 5'b01111; w[21][62] = 5'b10000; w[21][63] = 5'b00000; w[21][64] = 5'b01111; w[21][65] = 5'b00000; w[21][66] = 5'b00000; w[21][67] = 5'b01111; w[21][68] = 5'b01111; w[21][69] = 5'b01111; w[21][70] = 5'b01111; w[21][71] = 5'b01111; w[21][72] = 5'b01111; w[21][73] = 5'b00000; w[21][74] = 5'b01111; w[21][75] = 5'b01111; w[21][76] = 5'b10000; w[21][77] = 5'b00000; w[21][78] = 5'b01111; w[21][79] = 5'b01111; w[21][80] = 5'b00000; w[21][81] = 5'b01111; w[21][82] = 5'b01111; w[21][83] = 5'b01111; w[21][84] = 5'b01111; w[21][85] = 5'b01111; w[21][86] = 5'b01111; w[21][87] = 5'b00000; w[21][88] = 5'b01111; w[21][89] = 5'b01111; w[21][90] = 5'b10000; w[21][91] = 5'b10000; w[21][92] = 5'b01111; w[21][93] = 5'b01111; w[21][94] = 5'b01111; w[21][95] = 5'b01111; w[21][96] = 5'b01111; w[21][97] = 5'b01111; w[21][98] = 5'b01111; w[21][99] = 5'b01111; w[21][100] = 5'b01111; w[21][101] = 5'b00000; w[21][102] = 5'b01111; w[21][103] = 5'b01111; w[21][104] = 5'b10000; w[21][105] = 5'b10000; w[21][106] = 5'b01111; w[21][107] = 5'b00000; w[21][108] = 5'b00000; w[21][109] = 5'b01111; w[21][110] = 5'b01111; w[21][111] = 5'b01111; w[21][112] = 5'b01111; w[21][113] = 5'b01111; w[21][114] = 5'b01111; w[21][115] = 5'b00000; w[21][116] = 5'b01111; w[21][117] = 5'b01111; w[21][118] = 5'b10000; w[21][119] = 5'b10000; w[21][120] = 5'b00000; w[21][121] = 5'b00000; w[21][122] = 5'b00000; w[21][123] = 5'b01111; w[21][124] = 5'b01111; w[21][125] = 5'b01111; w[21][126] = 5'b01111; w[21][127] = 5'b01111; w[21][128] = 5'b01111; w[21][129] = 5'b00000; w[21][130] = 5'b01111; w[21][131] = 5'b01111; w[21][132] = 5'b00000; w[21][133] = 5'b10000; w[21][134] = 5'b01111; w[21][135] = 5'b01111; w[21][136] = 5'b00000; w[21][137] = 5'b01111; w[21][138] = 5'b01111; w[21][139] = 5'b01111; w[21][140] = 5'b01111; w[21][141] = 5'b01111; w[21][142] = 5'b01111; w[21][143] = 5'b00000; w[21][144] = 5'b00000; w[21][145] = 5'b01111; w[21][146] = 5'b00000; w[21][147] = 5'b10000; w[21][148] = 5'b01111; w[21][149] = 5'b00000; w[21][150] = 5'b00000; w[21][151] = 5'b01111; w[21][152] = 5'b01111; w[21][153] = 5'b01111; w[21][154] = 5'b01111; w[21][155] = 5'b01111; w[21][156] = 5'b01111; w[21][157] = 5'b00000; w[21][158] = 5'b00000; w[21][159] = 5'b00000; w[21][160] = 5'b10000; w[21][161] = 5'b10000; w[21][162] = 5'b10000; w[21][163] = 5'b00000; w[21][164] = 5'b00000; w[21][165] = 5'b01111; w[21][166] = 5'b01111; w[21][167] = 5'b01111; w[21][168] = 5'b01111; w[21][169] = 5'b01111; w[21][170] = 5'b01111; w[21][171] = 5'b01111; w[21][172] = 5'b00000; w[21][173] = 5'b00000; w[21][174] = 5'b10000; w[21][175] = 5'b10000; w[21][176] = 5'b10000; w[21][177] = 5'b00000; w[21][178] = 5'b01111; w[21][179] = 5'b01111; w[21][180] = 5'b01111; w[21][181] = 5'b01111; w[21][182] = 5'b01111; w[21][183] = 5'b01111; w[21][184] = 5'b01111; w[21][185] = 5'b01111; w[21][186] = 5'b01111; w[21][187] = 5'b01111; w[21][188] = 5'b01111; w[21][189] = 5'b01111; w[21][190] = 5'b01111; w[21][191] = 5'b01111; w[21][192] = 5'b01111; w[21][193] = 5'b01111; w[21][194] = 5'b01111; w[21][195] = 5'b01111; w[21][196] = 5'b01111; w[21][197] = 5'b01111; w[21][198] = 5'b01111; w[21][199] = 5'b01111; w[21][200] = 5'b01111; w[21][201] = 5'b01111; w[21][202] = 5'b01111; w[21][203] = 5'b01111; w[21][204] = 5'b01111; w[21][205] = 5'b01111; w[21][206] = 5'b01111; w[21][207] = 5'b01111; w[21][208] = 5'b01111; w[21][209] = 5'b01111; 
w[22][0] = 5'b01111; w[22][1] = 5'b01111; w[22][2] = 5'b01111; w[22][3] = 5'b01111; w[22][4] = 5'b01111; w[22][5] = 5'b01111; w[22][6] = 5'b01111; w[22][7] = 5'b01111; w[22][8] = 5'b01111; w[22][9] = 5'b01111; w[22][10] = 5'b01111; w[22][11] = 5'b01111; w[22][12] = 5'b01111; w[22][13] = 5'b01111; w[22][14] = 5'b01111; w[22][15] = 5'b01111; w[22][16] = 5'b01111; w[22][17] = 5'b01111; w[22][18] = 5'b01111; w[22][19] = 5'b01111; w[22][20] = 5'b01111; w[22][21] = 5'b01111; w[22][22] = 5'b00000; w[22][23] = 5'b01111; w[22][24] = 5'b01111; w[22][25] = 5'b01111; w[22][26] = 5'b01111; w[22][27] = 5'b01111; w[22][28] = 5'b01111; w[22][29] = 5'b01111; w[22][30] = 5'b01111; w[22][31] = 5'b00000; w[22][32] = 5'b10000; w[22][33] = 5'b10000; w[22][34] = 5'b10000; w[22][35] = 5'b10000; w[22][36] = 5'b10000; w[22][37] = 5'b10000; w[22][38] = 5'b00000; w[22][39] = 5'b01111; w[22][40] = 5'b01111; w[22][41] = 5'b01111; w[22][42] = 5'b01111; w[22][43] = 5'b01111; w[22][44] = 5'b01111; w[22][45] = 5'b10000; w[22][46] = 5'b10000; w[22][47] = 5'b10000; w[22][48] = 5'b10000; w[22][49] = 5'b10000; w[22][50] = 5'b10000; w[22][51] = 5'b10000; w[22][52] = 5'b10000; w[22][53] = 5'b01111; w[22][54] = 5'b01111; w[22][55] = 5'b01111; w[22][56] = 5'b01111; w[22][57] = 5'b01111; w[22][58] = 5'b01111; w[22][59] = 5'b00000; w[22][60] = 5'b00000; w[22][61] = 5'b01111; w[22][62] = 5'b10000; w[22][63] = 5'b00000; w[22][64] = 5'b01111; w[22][65] = 5'b00000; w[22][66] = 5'b00000; w[22][67] = 5'b01111; w[22][68] = 5'b01111; w[22][69] = 5'b01111; w[22][70] = 5'b01111; w[22][71] = 5'b01111; w[22][72] = 5'b01111; w[22][73] = 5'b00000; w[22][74] = 5'b01111; w[22][75] = 5'b01111; w[22][76] = 5'b10000; w[22][77] = 5'b00000; w[22][78] = 5'b01111; w[22][79] = 5'b01111; w[22][80] = 5'b00000; w[22][81] = 5'b01111; w[22][82] = 5'b01111; w[22][83] = 5'b01111; w[22][84] = 5'b01111; w[22][85] = 5'b01111; w[22][86] = 5'b01111; w[22][87] = 5'b00000; w[22][88] = 5'b01111; w[22][89] = 5'b01111; w[22][90] = 5'b10000; w[22][91] = 5'b10000; w[22][92] = 5'b01111; w[22][93] = 5'b01111; w[22][94] = 5'b01111; w[22][95] = 5'b01111; w[22][96] = 5'b01111; w[22][97] = 5'b01111; w[22][98] = 5'b01111; w[22][99] = 5'b01111; w[22][100] = 5'b01111; w[22][101] = 5'b00000; w[22][102] = 5'b01111; w[22][103] = 5'b01111; w[22][104] = 5'b10000; w[22][105] = 5'b10000; w[22][106] = 5'b01111; w[22][107] = 5'b00000; w[22][108] = 5'b00000; w[22][109] = 5'b01111; w[22][110] = 5'b01111; w[22][111] = 5'b01111; w[22][112] = 5'b01111; w[22][113] = 5'b01111; w[22][114] = 5'b01111; w[22][115] = 5'b00000; w[22][116] = 5'b01111; w[22][117] = 5'b01111; w[22][118] = 5'b10000; w[22][119] = 5'b10000; w[22][120] = 5'b00000; w[22][121] = 5'b00000; w[22][122] = 5'b00000; w[22][123] = 5'b01111; w[22][124] = 5'b01111; w[22][125] = 5'b01111; w[22][126] = 5'b01111; w[22][127] = 5'b01111; w[22][128] = 5'b01111; w[22][129] = 5'b00000; w[22][130] = 5'b01111; w[22][131] = 5'b01111; w[22][132] = 5'b00000; w[22][133] = 5'b10000; w[22][134] = 5'b01111; w[22][135] = 5'b01111; w[22][136] = 5'b00000; w[22][137] = 5'b01111; w[22][138] = 5'b01111; w[22][139] = 5'b01111; w[22][140] = 5'b01111; w[22][141] = 5'b01111; w[22][142] = 5'b01111; w[22][143] = 5'b00000; w[22][144] = 5'b00000; w[22][145] = 5'b01111; w[22][146] = 5'b00000; w[22][147] = 5'b10000; w[22][148] = 5'b01111; w[22][149] = 5'b00000; w[22][150] = 5'b00000; w[22][151] = 5'b01111; w[22][152] = 5'b01111; w[22][153] = 5'b01111; w[22][154] = 5'b01111; w[22][155] = 5'b01111; w[22][156] = 5'b01111; w[22][157] = 5'b00000; w[22][158] = 5'b00000; w[22][159] = 5'b00000; w[22][160] = 5'b10000; w[22][161] = 5'b10000; w[22][162] = 5'b10000; w[22][163] = 5'b00000; w[22][164] = 5'b00000; w[22][165] = 5'b01111; w[22][166] = 5'b01111; w[22][167] = 5'b01111; w[22][168] = 5'b01111; w[22][169] = 5'b01111; w[22][170] = 5'b01111; w[22][171] = 5'b01111; w[22][172] = 5'b00000; w[22][173] = 5'b00000; w[22][174] = 5'b10000; w[22][175] = 5'b10000; w[22][176] = 5'b10000; w[22][177] = 5'b00000; w[22][178] = 5'b01111; w[22][179] = 5'b01111; w[22][180] = 5'b01111; w[22][181] = 5'b01111; w[22][182] = 5'b01111; w[22][183] = 5'b01111; w[22][184] = 5'b01111; w[22][185] = 5'b01111; w[22][186] = 5'b01111; w[22][187] = 5'b01111; w[22][188] = 5'b01111; w[22][189] = 5'b01111; w[22][190] = 5'b01111; w[22][191] = 5'b01111; w[22][192] = 5'b01111; w[22][193] = 5'b01111; w[22][194] = 5'b01111; w[22][195] = 5'b01111; w[22][196] = 5'b01111; w[22][197] = 5'b01111; w[22][198] = 5'b01111; w[22][199] = 5'b01111; w[22][200] = 5'b01111; w[22][201] = 5'b01111; w[22][202] = 5'b01111; w[22][203] = 5'b01111; w[22][204] = 5'b01111; w[22][205] = 5'b01111; w[22][206] = 5'b01111; w[22][207] = 5'b01111; w[22][208] = 5'b01111; w[22][209] = 5'b01111; 
w[23][0] = 5'b01111; w[23][1] = 5'b01111; w[23][2] = 5'b01111; w[23][3] = 5'b01111; w[23][4] = 5'b01111; w[23][5] = 5'b01111; w[23][6] = 5'b01111; w[23][7] = 5'b01111; w[23][8] = 5'b01111; w[23][9] = 5'b01111; w[23][10] = 5'b01111; w[23][11] = 5'b01111; w[23][12] = 5'b01111; w[23][13] = 5'b01111; w[23][14] = 5'b01111; w[23][15] = 5'b01111; w[23][16] = 5'b01111; w[23][17] = 5'b01111; w[23][18] = 5'b01111; w[23][19] = 5'b01111; w[23][20] = 5'b01111; w[23][21] = 5'b01111; w[23][22] = 5'b01111; w[23][23] = 5'b00000; w[23][24] = 5'b01111; w[23][25] = 5'b01111; w[23][26] = 5'b01111; w[23][27] = 5'b01111; w[23][28] = 5'b01111; w[23][29] = 5'b01111; w[23][30] = 5'b01111; w[23][31] = 5'b00000; w[23][32] = 5'b10000; w[23][33] = 5'b10000; w[23][34] = 5'b10000; w[23][35] = 5'b10000; w[23][36] = 5'b10000; w[23][37] = 5'b10000; w[23][38] = 5'b00000; w[23][39] = 5'b01111; w[23][40] = 5'b01111; w[23][41] = 5'b01111; w[23][42] = 5'b01111; w[23][43] = 5'b01111; w[23][44] = 5'b01111; w[23][45] = 5'b10000; w[23][46] = 5'b10000; w[23][47] = 5'b10000; w[23][48] = 5'b10000; w[23][49] = 5'b10000; w[23][50] = 5'b10000; w[23][51] = 5'b10000; w[23][52] = 5'b10000; w[23][53] = 5'b01111; w[23][54] = 5'b01111; w[23][55] = 5'b01111; w[23][56] = 5'b01111; w[23][57] = 5'b01111; w[23][58] = 5'b01111; w[23][59] = 5'b00000; w[23][60] = 5'b00000; w[23][61] = 5'b01111; w[23][62] = 5'b10000; w[23][63] = 5'b00000; w[23][64] = 5'b01111; w[23][65] = 5'b00000; w[23][66] = 5'b00000; w[23][67] = 5'b01111; w[23][68] = 5'b01111; w[23][69] = 5'b01111; w[23][70] = 5'b01111; w[23][71] = 5'b01111; w[23][72] = 5'b01111; w[23][73] = 5'b00000; w[23][74] = 5'b01111; w[23][75] = 5'b01111; w[23][76] = 5'b10000; w[23][77] = 5'b00000; w[23][78] = 5'b01111; w[23][79] = 5'b01111; w[23][80] = 5'b00000; w[23][81] = 5'b01111; w[23][82] = 5'b01111; w[23][83] = 5'b01111; w[23][84] = 5'b01111; w[23][85] = 5'b01111; w[23][86] = 5'b01111; w[23][87] = 5'b00000; w[23][88] = 5'b01111; w[23][89] = 5'b01111; w[23][90] = 5'b10000; w[23][91] = 5'b10000; w[23][92] = 5'b01111; w[23][93] = 5'b01111; w[23][94] = 5'b01111; w[23][95] = 5'b01111; w[23][96] = 5'b01111; w[23][97] = 5'b01111; w[23][98] = 5'b01111; w[23][99] = 5'b01111; w[23][100] = 5'b01111; w[23][101] = 5'b00000; w[23][102] = 5'b01111; w[23][103] = 5'b01111; w[23][104] = 5'b10000; w[23][105] = 5'b10000; w[23][106] = 5'b01111; w[23][107] = 5'b00000; w[23][108] = 5'b00000; w[23][109] = 5'b01111; w[23][110] = 5'b01111; w[23][111] = 5'b01111; w[23][112] = 5'b01111; w[23][113] = 5'b01111; w[23][114] = 5'b01111; w[23][115] = 5'b00000; w[23][116] = 5'b01111; w[23][117] = 5'b01111; w[23][118] = 5'b10000; w[23][119] = 5'b10000; w[23][120] = 5'b00000; w[23][121] = 5'b00000; w[23][122] = 5'b00000; w[23][123] = 5'b01111; w[23][124] = 5'b01111; w[23][125] = 5'b01111; w[23][126] = 5'b01111; w[23][127] = 5'b01111; w[23][128] = 5'b01111; w[23][129] = 5'b00000; w[23][130] = 5'b01111; w[23][131] = 5'b01111; w[23][132] = 5'b00000; w[23][133] = 5'b10000; w[23][134] = 5'b01111; w[23][135] = 5'b01111; w[23][136] = 5'b00000; w[23][137] = 5'b01111; w[23][138] = 5'b01111; w[23][139] = 5'b01111; w[23][140] = 5'b01111; w[23][141] = 5'b01111; w[23][142] = 5'b01111; w[23][143] = 5'b00000; w[23][144] = 5'b00000; w[23][145] = 5'b01111; w[23][146] = 5'b00000; w[23][147] = 5'b10000; w[23][148] = 5'b01111; w[23][149] = 5'b00000; w[23][150] = 5'b00000; w[23][151] = 5'b01111; w[23][152] = 5'b01111; w[23][153] = 5'b01111; w[23][154] = 5'b01111; w[23][155] = 5'b01111; w[23][156] = 5'b01111; w[23][157] = 5'b00000; w[23][158] = 5'b00000; w[23][159] = 5'b00000; w[23][160] = 5'b10000; w[23][161] = 5'b10000; w[23][162] = 5'b10000; w[23][163] = 5'b00000; w[23][164] = 5'b00000; w[23][165] = 5'b01111; w[23][166] = 5'b01111; w[23][167] = 5'b01111; w[23][168] = 5'b01111; w[23][169] = 5'b01111; w[23][170] = 5'b01111; w[23][171] = 5'b01111; w[23][172] = 5'b00000; w[23][173] = 5'b00000; w[23][174] = 5'b10000; w[23][175] = 5'b10000; w[23][176] = 5'b10000; w[23][177] = 5'b00000; w[23][178] = 5'b01111; w[23][179] = 5'b01111; w[23][180] = 5'b01111; w[23][181] = 5'b01111; w[23][182] = 5'b01111; w[23][183] = 5'b01111; w[23][184] = 5'b01111; w[23][185] = 5'b01111; w[23][186] = 5'b01111; w[23][187] = 5'b01111; w[23][188] = 5'b01111; w[23][189] = 5'b01111; w[23][190] = 5'b01111; w[23][191] = 5'b01111; w[23][192] = 5'b01111; w[23][193] = 5'b01111; w[23][194] = 5'b01111; w[23][195] = 5'b01111; w[23][196] = 5'b01111; w[23][197] = 5'b01111; w[23][198] = 5'b01111; w[23][199] = 5'b01111; w[23][200] = 5'b01111; w[23][201] = 5'b01111; w[23][202] = 5'b01111; w[23][203] = 5'b01111; w[23][204] = 5'b01111; w[23][205] = 5'b01111; w[23][206] = 5'b01111; w[23][207] = 5'b01111; w[23][208] = 5'b01111; w[23][209] = 5'b01111; 
w[24][0] = 5'b01111; w[24][1] = 5'b01111; w[24][2] = 5'b01111; w[24][3] = 5'b01111; w[24][4] = 5'b01111; w[24][5] = 5'b01111; w[24][6] = 5'b01111; w[24][7] = 5'b01111; w[24][8] = 5'b01111; w[24][9] = 5'b01111; w[24][10] = 5'b01111; w[24][11] = 5'b01111; w[24][12] = 5'b01111; w[24][13] = 5'b01111; w[24][14] = 5'b01111; w[24][15] = 5'b01111; w[24][16] = 5'b01111; w[24][17] = 5'b01111; w[24][18] = 5'b01111; w[24][19] = 5'b01111; w[24][20] = 5'b01111; w[24][21] = 5'b01111; w[24][22] = 5'b01111; w[24][23] = 5'b01111; w[24][24] = 5'b00000; w[24][25] = 5'b01111; w[24][26] = 5'b01111; w[24][27] = 5'b01111; w[24][28] = 5'b01111; w[24][29] = 5'b01111; w[24][30] = 5'b01111; w[24][31] = 5'b00000; w[24][32] = 5'b10000; w[24][33] = 5'b10000; w[24][34] = 5'b10000; w[24][35] = 5'b10000; w[24][36] = 5'b10000; w[24][37] = 5'b10000; w[24][38] = 5'b00000; w[24][39] = 5'b01111; w[24][40] = 5'b01111; w[24][41] = 5'b01111; w[24][42] = 5'b01111; w[24][43] = 5'b01111; w[24][44] = 5'b01111; w[24][45] = 5'b10000; w[24][46] = 5'b10000; w[24][47] = 5'b10000; w[24][48] = 5'b10000; w[24][49] = 5'b10000; w[24][50] = 5'b10000; w[24][51] = 5'b10000; w[24][52] = 5'b10000; w[24][53] = 5'b01111; w[24][54] = 5'b01111; w[24][55] = 5'b01111; w[24][56] = 5'b01111; w[24][57] = 5'b01111; w[24][58] = 5'b01111; w[24][59] = 5'b00000; w[24][60] = 5'b00000; w[24][61] = 5'b01111; w[24][62] = 5'b10000; w[24][63] = 5'b00000; w[24][64] = 5'b01111; w[24][65] = 5'b00000; w[24][66] = 5'b00000; w[24][67] = 5'b01111; w[24][68] = 5'b01111; w[24][69] = 5'b01111; w[24][70] = 5'b01111; w[24][71] = 5'b01111; w[24][72] = 5'b01111; w[24][73] = 5'b00000; w[24][74] = 5'b01111; w[24][75] = 5'b01111; w[24][76] = 5'b10000; w[24][77] = 5'b00000; w[24][78] = 5'b01111; w[24][79] = 5'b01111; w[24][80] = 5'b00000; w[24][81] = 5'b01111; w[24][82] = 5'b01111; w[24][83] = 5'b01111; w[24][84] = 5'b01111; w[24][85] = 5'b01111; w[24][86] = 5'b01111; w[24][87] = 5'b00000; w[24][88] = 5'b01111; w[24][89] = 5'b01111; w[24][90] = 5'b10000; w[24][91] = 5'b10000; w[24][92] = 5'b01111; w[24][93] = 5'b01111; w[24][94] = 5'b01111; w[24][95] = 5'b01111; w[24][96] = 5'b01111; w[24][97] = 5'b01111; w[24][98] = 5'b01111; w[24][99] = 5'b01111; w[24][100] = 5'b01111; w[24][101] = 5'b00000; w[24][102] = 5'b01111; w[24][103] = 5'b01111; w[24][104] = 5'b10000; w[24][105] = 5'b10000; w[24][106] = 5'b01111; w[24][107] = 5'b00000; w[24][108] = 5'b00000; w[24][109] = 5'b01111; w[24][110] = 5'b01111; w[24][111] = 5'b01111; w[24][112] = 5'b01111; w[24][113] = 5'b01111; w[24][114] = 5'b01111; w[24][115] = 5'b00000; w[24][116] = 5'b01111; w[24][117] = 5'b01111; w[24][118] = 5'b10000; w[24][119] = 5'b10000; w[24][120] = 5'b00000; w[24][121] = 5'b00000; w[24][122] = 5'b00000; w[24][123] = 5'b01111; w[24][124] = 5'b01111; w[24][125] = 5'b01111; w[24][126] = 5'b01111; w[24][127] = 5'b01111; w[24][128] = 5'b01111; w[24][129] = 5'b00000; w[24][130] = 5'b01111; w[24][131] = 5'b01111; w[24][132] = 5'b00000; w[24][133] = 5'b10000; w[24][134] = 5'b01111; w[24][135] = 5'b01111; w[24][136] = 5'b00000; w[24][137] = 5'b01111; w[24][138] = 5'b01111; w[24][139] = 5'b01111; w[24][140] = 5'b01111; w[24][141] = 5'b01111; w[24][142] = 5'b01111; w[24][143] = 5'b00000; w[24][144] = 5'b00000; w[24][145] = 5'b01111; w[24][146] = 5'b00000; w[24][147] = 5'b10000; w[24][148] = 5'b01111; w[24][149] = 5'b00000; w[24][150] = 5'b00000; w[24][151] = 5'b01111; w[24][152] = 5'b01111; w[24][153] = 5'b01111; w[24][154] = 5'b01111; w[24][155] = 5'b01111; w[24][156] = 5'b01111; w[24][157] = 5'b00000; w[24][158] = 5'b00000; w[24][159] = 5'b00000; w[24][160] = 5'b10000; w[24][161] = 5'b10000; w[24][162] = 5'b10000; w[24][163] = 5'b00000; w[24][164] = 5'b00000; w[24][165] = 5'b01111; w[24][166] = 5'b01111; w[24][167] = 5'b01111; w[24][168] = 5'b01111; w[24][169] = 5'b01111; w[24][170] = 5'b01111; w[24][171] = 5'b01111; w[24][172] = 5'b00000; w[24][173] = 5'b00000; w[24][174] = 5'b10000; w[24][175] = 5'b10000; w[24][176] = 5'b10000; w[24][177] = 5'b00000; w[24][178] = 5'b01111; w[24][179] = 5'b01111; w[24][180] = 5'b01111; w[24][181] = 5'b01111; w[24][182] = 5'b01111; w[24][183] = 5'b01111; w[24][184] = 5'b01111; w[24][185] = 5'b01111; w[24][186] = 5'b01111; w[24][187] = 5'b01111; w[24][188] = 5'b01111; w[24][189] = 5'b01111; w[24][190] = 5'b01111; w[24][191] = 5'b01111; w[24][192] = 5'b01111; w[24][193] = 5'b01111; w[24][194] = 5'b01111; w[24][195] = 5'b01111; w[24][196] = 5'b01111; w[24][197] = 5'b01111; w[24][198] = 5'b01111; w[24][199] = 5'b01111; w[24][200] = 5'b01111; w[24][201] = 5'b01111; w[24][202] = 5'b01111; w[24][203] = 5'b01111; w[24][204] = 5'b01111; w[24][205] = 5'b01111; w[24][206] = 5'b01111; w[24][207] = 5'b01111; w[24][208] = 5'b01111; w[24][209] = 5'b01111; 
w[25][0] = 5'b01111; w[25][1] = 5'b01111; w[25][2] = 5'b01111; w[25][3] = 5'b01111; w[25][4] = 5'b01111; w[25][5] = 5'b01111; w[25][6] = 5'b01111; w[25][7] = 5'b01111; w[25][8] = 5'b01111; w[25][9] = 5'b01111; w[25][10] = 5'b01111; w[25][11] = 5'b01111; w[25][12] = 5'b01111; w[25][13] = 5'b01111; w[25][14] = 5'b01111; w[25][15] = 5'b01111; w[25][16] = 5'b01111; w[25][17] = 5'b01111; w[25][18] = 5'b01111; w[25][19] = 5'b01111; w[25][20] = 5'b01111; w[25][21] = 5'b01111; w[25][22] = 5'b01111; w[25][23] = 5'b01111; w[25][24] = 5'b01111; w[25][25] = 5'b00000; w[25][26] = 5'b01111; w[25][27] = 5'b01111; w[25][28] = 5'b01111; w[25][29] = 5'b01111; w[25][30] = 5'b01111; w[25][31] = 5'b00000; w[25][32] = 5'b10000; w[25][33] = 5'b10000; w[25][34] = 5'b10000; w[25][35] = 5'b10000; w[25][36] = 5'b10000; w[25][37] = 5'b10000; w[25][38] = 5'b00000; w[25][39] = 5'b01111; w[25][40] = 5'b01111; w[25][41] = 5'b01111; w[25][42] = 5'b01111; w[25][43] = 5'b01111; w[25][44] = 5'b01111; w[25][45] = 5'b10000; w[25][46] = 5'b10000; w[25][47] = 5'b10000; w[25][48] = 5'b10000; w[25][49] = 5'b10000; w[25][50] = 5'b10000; w[25][51] = 5'b10000; w[25][52] = 5'b10000; w[25][53] = 5'b01111; w[25][54] = 5'b01111; w[25][55] = 5'b01111; w[25][56] = 5'b01111; w[25][57] = 5'b01111; w[25][58] = 5'b01111; w[25][59] = 5'b00000; w[25][60] = 5'b00000; w[25][61] = 5'b01111; w[25][62] = 5'b10000; w[25][63] = 5'b00000; w[25][64] = 5'b01111; w[25][65] = 5'b00000; w[25][66] = 5'b00000; w[25][67] = 5'b01111; w[25][68] = 5'b01111; w[25][69] = 5'b01111; w[25][70] = 5'b01111; w[25][71] = 5'b01111; w[25][72] = 5'b01111; w[25][73] = 5'b00000; w[25][74] = 5'b01111; w[25][75] = 5'b01111; w[25][76] = 5'b10000; w[25][77] = 5'b00000; w[25][78] = 5'b01111; w[25][79] = 5'b01111; w[25][80] = 5'b00000; w[25][81] = 5'b01111; w[25][82] = 5'b01111; w[25][83] = 5'b01111; w[25][84] = 5'b01111; w[25][85] = 5'b01111; w[25][86] = 5'b01111; w[25][87] = 5'b00000; w[25][88] = 5'b01111; w[25][89] = 5'b01111; w[25][90] = 5'b10000; w[25][91] = 5'b10000; w[25][92] = 5'b01111; w[25][93] = 5'b01111; w[25][94] = 5'b01111; w[25][95] = 5'b01111; w[25][96] = 5'b01111; w[25][97] = 5'b01111; w[25][98] = 5'b01111; w[25][99] = 5'b01111; w[25][100] = 5'b01111; w[25][101] = 5'b00000; w[25][102] = 5'b01111; w[25][103] = 5'b01111; w[25][104] = 5'b10000; w[25][105] = 5'b10000; w[25][106] = 5'b01111; w[25][107] = 5'b00000; w[25][108] = 5'b00000; w[25][109] = 5'b01111; w[25][110] = 5'b01111; w[25][111] = 5'b01111; w[25][112] = 5'b01111; w[25][113] = 5'b01111; w[25][114] = 5'b01111; w[25][115] = 5'b00000; w[25][116] = 5'b01111; w[25][117] = 5'b01111; w[25][118] = 5'b10000; w[25][119] = 5'b10000; w[25][120] = 5'b00000; w[25][121] = 5'b00000; w[25][122] = 5'b00000; w[25][123] = 5'b01111; w[25][124] = 5'b01111; w[25][125] = 5'b01111; w[25][126] = 5'b01111; w[25][127] = 5'b01111; w[25][128] = 5'b01111; w[25][129] = 5'b00000; w[25][130] = 5'b01111; w[25][131] = 5'b01111; w[25][132] = 5'b00000; w[25][133] = 5'b10000; w[25][134] = 5'b01111; w[25][135] = 5'b01111; w[25][136] = 5'b00000; w[25][137] = 5'b01111; w[25][138] = 5'b01111; w[25][139] = 5'b01111; w[25][140] = 5'b01111; w[25][141] = 5'b01111; w[25][142] = 5'b01111; w[25][143] = 5'b00000; w[25][144] = 5'b00000; w[25][145] = 5'b01111; w[25][146] = 5'b00000; w[25][147] = 5'b10000; w[25][148] = 5'b01111; w[25][149] = 5'b00000; w[25][150] = 5'b00000; w[25][151] = 5'b01111; w[25][152] = 5'b01111; w[25][153] = 5'b01111; w[25][154] = 5'b01111; w[25][155] = 5'b01111; w[25][156] = 5'b01111; w[25][157] = 5'b00000; w[25][158] = 5'b00000; w[25][159] = 5'b00000; w[25][160] = 5'b10000; w[25][161] = 5'b10000; w[25][162] = 5'b10000; w[25][163] = 5'b00000; w[25][164] = 5'b00000; w[25][165] = 5'b01111; w[25][166] = 5'b01111; w[25][167] = 5'b01111; w[25][168] = 5'b01111; w[25][169] = 5'b01111; w[25][170] = 5'b01111; w[25][171] = 5'b01111; w[25][172] = 5'b00000; w[25][173] = 5'b00000; w[25][174] = 5'b10000; w[25][175] = 5'b10000; w[25][176] = 5'b10000; w[25][177] = 5'b00000; w[25][178] = 5'b01111; w[25][179] = 5'b01111; w[25][180] = 5'b01111; w[25][181] = 5'b01111; w[25][182] = 5'b01111; w[25][183] = 5'b01111; w[25][184] = 5'b01111; w[25][185] = 5'b01111; w[25][186] = 5'b01111; w[25][187] = 5'b01111; w[25][188] = 5'b01111; w[25][189] = 5'b01111; w[25][190] = 5'b01111; w[25][191] = 5'b01111; w[25][192] = 5'b01111; w[25][193] = 5'b01111; w[25][194] = 5'b01111; w[25][195] = 5'b01111; w[25][196] = 5'b01111; w[25][197] = 5'b01111; w[25][198] = 5'b01111; w[25][199] = 5'b01111; w[25][200] = 5'b01111; w[25][201] = 5'b01111; w[25][202] = 5'b01111; w[25][203] = 5'b01111; w[25][204] = 5'b01111; w[25][205] = 5'b01111; w[25][206] = 5'b01111; w[25][207] = 5'b01111; w[25][208] = 5'b01111; w[25][209] = 5'b01111; 
w[26][0] = 5'b01111; w[26][1] = 5'b01111; w[26][2] = 5'b01111; w[26][3] = 5'b01111; w[26][4] = 5'b01111; w[26][5] = 5'b01111; w[26][6] = 5'b01111; w[26][7] = 5'b01111; w[26][8] = 5'b01111; w[26][9] = 5'b01111; w[26][10] = 5'b01111; w[26][11] = 5'b01111; w[26][12] = 5'b01111; w[26][13] = 5'b01111; w[26][14] = 5'b01111; w[26][15] = 5'b01111; w[26][16] = 5'b01111; w[26][17] = 5'b01111; w[26][18] = 5'b01111; w[26][19] = 5'b01111; w[26][20] = 5'b01111; w[26][21] = 5'b01111; w[26][22] = 5'b01111; w[26][23] = 5'b01111; w[26][24] = 5'b01111; w[26][25] = 5'b01111; w[26][26] = 5'b00000; w[26][27] = 5'b01111; w[26][28] = 5'b01111; w[26][29] = 5'b01111; w[26][30] = 5'b01111; w[26][31] = 5'b00000; w[26][32] = 5'b10000; w[26][33] = 5'b10000; w[26][34] = 5'b10000; w[26][35] = 5'b10000; w[26][36] = 5'b10000; w[26][37] = 5'b10000; w[26][38] = 5'b00000; w[26][39] = 5'b01111; w[26][40] = 5'b01111; w[26][41] = 5'b01111; w[26][42] = 5'b01111; w[26][43] = 5'b01111; w[26][44] = 5'b01111; w[26][45] = 5'b10000; w[26][46] = 5'b10000; w[26][47] = 5'b10000; w[26][48] = 5'b10000; w[26][49] = 5'b10000; w[26][50] = 5'b10000; w[26][51] = 5'b10000; w[26][52] = 5'b10000; w[26][53] = 5'b01111; w[26][54] = 5'b01111; w[26][55] = 5'b01111; w[26][56] = 5'b01111; w[26][57] = 5'b01111; w[26][58] = 5'b01111; w[26][59] = 5'b00000; w[26][60] = 5'b00000; w[26][61] = 5'b01111; w[26][62] = 5'b10000; w[26][63] = 5'b00000; w[26][64] = 5'b01111; w[26][65] = 5'b00000; w[26][66] = 5'b00000; w[26][67] = 5'b01111; w[26][68] = 5'b01111; w[26][69] = 5'b01111; w[26][70] = 5'b01111; w[26][71] = 5'b01111; w[26][72] = 5'b01111; w[26][73] = 5'b00000; w[26][74] = 5'b01111; w[26][75] = 5'b01111; w[26][76] = 5'b10000; w[26][77] = 5'b00000; w[26][78] = 5'b01111; w[26][79] = 5'b01111; w[26][80] = 5'b00000; w[26][81] = 5'b01111; w[26][82] = 5'b01111; w[26][83] = 5'b01111; w[26][84] = 5'b01111; w[26][85] = 5'b01111; w[26][86] = 5'b01111; w[26][87] = 5'b00000; w[26][88] = 5'b01111; w[26][89] = 5'b01111; w[26][90] = 5'b10000; w[26][91] = 5'b10000; w[26][92] = 5'b01111; w[26][93] = 5'b01111; w[26][94] = 5'b01111; w[26][95] = 5'b01111; w[26][96] = 5'b01111; w[26][97] = 5'b01111; w[26][98] = 5'b01111; w[26][99] = 5'b01111; w[26][100] = 5'b01111; w[26][101] = 5'b00000; w[26][102] = 5'b01111; w[26][103] = 5'b01111; w[26][104] = 5'b10000; w[26][105] = 5'b10000; w[26][106] = 5'b01111; w[26][107] = 5'b00000; w[26][108] = 5'b00000; w[26][109] = 5'b01111; w[26][110] = 5'b01111; w[26][111] = 5'b01111; w[26][112] = 5'b01111; w[26][113] = 5'b01111; w[26][114] = 5'b01111; w[26][115] = 5'b00000; w[26][116] = 5'b01111; w[26][117] = 5'b01111; w[26][118] = 5'b10000; w[26][119] = 5'b10000; w[26][120] = 5'b00000; w[26][121] = 5'b00000; w[26][122] = 5'b00000; w[26][123] = 5'b01111; w[26][124] = 5'b01111; w[26][125] = 5'b01111; w[26][126] = 5'b01111; w[26][127] = 5'b01111; w[26][128] = 5'b01111; w[26][129] = 5'b00000; w[26][130] = 5'b01111; w[26][131] = 5'b01111; w[26][132] = 5'b00000; w[26][133] = 5'b10000; w[26][134] = 5'b01111; w[26][135] = 5'b01111; w[26][136] = 5'b00000; w[26][137] = 5'b01111; w[26][138] = 5'b01111; w[26][139] = 5'b01111; w[26][140] = 5'b01111; w[26][141] = 5'b01111; w[26][142] = 5'b01111; w[26][143] = 5'b00000; w[26][144] = 5'b00000; w[26][145] = 5'b01111; w[26][146] = 5'b00000; w[26][147] = 5'b10000; w[26][148] = 5'b01111; w[26][149] = 5'b00000; w[26][150] = 5'b00000; w[26][151] = 5'b01111; w[26][152] = 5'b01111; w[26][153] = 5'b01111; w[26][154] = 5'b01111; w[26][155] = 5'b01111; w[26][156] = 5'b01111; w[26][157] = 5'b00000; w[26][158] = 5'b00000; w[26][159] = 5'b00000; w[26][160] = 5'b10000; w[26][161] = 5'b10000; w[26][162] = 5'b10000; w[26][163] = 5'b00000; w[26][164] = 5'b00000; w[26][165] = 5'b01111; w[26][166] = 5'b01111; w[26][167] = 5'b01111; w[26][168] = 5'b01111; w[26][169] = 5'b01111; w[26][170] = 5'b01111; w[26][171] = 5'b01111; w[26][172] = 5'b00000; w[26][173] = 5'b00000; w[26][174] = 5'b10000; w[26][175] = 5'b10000; w[26][176] = 5'b10000; w[26][177] = 5'b00000; w[26][178] = 5'b01111; w[26][179] = 5'b01111; w[26][180] = 5'b01111; w[26][181] = 5'b01111; w[26][182] = 5'b01111; w[26][183] = 5'b01111; w[26][184] = 5'b01111; w[26][185] = 5'b01111; w[26][186] = 5'b01111; w[26][187] = 5'b01111; w[26][188] = 5'b01111; w[26][189] = 5'b01111; w[26][190] = 5'b01111; w[26][191] = 5'b01111; w[26][192] = 5'b01111; w[26][193] = 5'b01111; w[26][194] = 5'b01111; w[26][195] = 5'b01111; w[26][196] = 5'b01111; w[26][197] = 5'b01111; w[26][198] = 5'b01111; w[26][199] = 5'b01111; w[26][200] = 5'b01111; w[26][201] = 5'b01111; w[26][202] = 5'b01111; w[26][203] = 5'b01111; w[26][204] = 5'b01111; w[26][205] = 5'b01111; w[26][206] = 5'b01111; w[26][207] = 5'b01111; w[26][208] = 5'b01111; w[26][209] = 5'b01111; 
w[27][0] = 5'b01111; w[27][1] = 5'b01111; w[27][2] = 5'b01111; w[27][3] = 5'b01111; w[27][4] = 5'b01111; w[27][5] = 5'b01111; w[27][6] = 5'b01111; w[27][7] = 5'b01111; w[27][8] = 5'b01111; w[27][9] = 5'b01111; w[27][10] = 5'b01111; w[27][11] = 5'b01111; w[27][12] = 5'b01111; w[27][13] = 5'b01111; w[27][14] = 5'b01111; w[27][15] = 5'b01111; w[27][16] = 5'b01111; w[27][17] = 5'b01111; w[27][18] = 5'b01111; w[27][19] = 5'b01111; w[27][20] = 5'b01111; w[27][21] = 5'b01111; w[27][22] = 5'b01111; w[27][23] = 5'b01111; w[27][24] = 5'b01111; w[27][25] = 5'b01111; w[27][26] = 5'b01111; w[27][27] = 5'b00000; w[27][28] = 5'b01111; w[27][29] = 5'b01111; w[27][30] = 5'b01111; w[27][31] = 5'b00000; w[27][32] = 5'b10000; w[27][33] = 5'b10000; w[27][34] = 5'b10000; w[27][35] = 5'b10000; w[27][36] = 5'b10000; w[27][37] = 5'b10000; w[27][38] = 5'b00000; w[27][39] = 5'b01111; w[27][40] = 5'b01111; w[27][41] = 5'b01111; w[27][42] = 5'b01111; w[27][43] = 5'b01111; w[27][44] = 5'b01111; w[27][45] = 5'b10000; w[27][46] = 5'b10000; w[27][47] = 5'b10000; w[27][48] = 5'b10000; w[27][49] = 5'b10000; w[27][50] = 5'b10000; w[27][51] = 5'b10000; w[27][52] = 5'b10000; w[27][53] = 5'b01111; w[27][54] = 5'b01111; w[27][55] = 5'b01111; w[27][56] = 5'b01111; w[27][57] = 5'b01111; w[27][58] = 5'b01111; w[27][59] = 5'b00000; w[27][60] = 5'b00000; w[27][61] = 5'b01111; w[27][62] = 5'b10000; w[27][63] = 5'b00000; w[27][64] = 5'b01111; w[27][65] = 5'b00000; w[27][66] = 5'b00000; w[27][67] = 5'b01111; w[27][68] = 5'b01111; w[27][69] = 5'b01111; w[27][70] = 5'b01111; w[27][71] = 5'b01111; w[27][72] = 5'b01111; w[27][73] = 5'b00000; w[27][74] = 5'b01111; w[27][75] = 5'b01111; w[27][76] = 5'b10000; w[27][77] = 5'b00000; w[27][78] = 5'b01111; w[27][79] = 5'b01111; w[27][80] = 5'b00000; w[27][81] = 5'b01111; w[27][82] = 5'b01111; w[27][83] = 5'b01111; w[27][84] = 5'b01111; w[27][85] = 5'b01111; w[27][86] = 5'b01111; w[27][87] = 5'b00000; w[27][88] = 5'b01111; w[27][89] = 5'b01111; w[27][90] = 5'b10000; w[27][91] = 5'b10000; w[27][92] = 5'b01111; w[27][93] = 5'b01111; w[27][94] = 5'b01111; w[27][95] = 5'b01111; w[27][96] = 5'b01111; w[27][97] = 5'b01111; w[27][98] = 5'b01111; w[27][99] = 5'b01111; w[27][100] = 5'b01111; w[27][101] = 5'b00000; w[27][102] = 5'b01111; w[27][103] = 5'b01111; w[27][104] = 5'b10000; w[27][105] = 5'b10000; w[27][106] = 5'b01111; w[27][107] = 5'b00000; w[27][108] = 5'b00000; w[27][109] = 5'b01111; w[27][110] = 5'b01111; w[27][111] = 5'b01111; w[27][112] = 5'b01111; w[27][113] = 5'b01111; w[27][114] = 5'b01111; w[27][115] = 5'b00000; w[27][116] = 5'b01111; w[27][117] = 5'b01111; w[27][118] = 5'b10000; w[27][119] = 5'b10000; w[27][120] = 5'b00000; w[27][121] = 5'b00000; w[27][122] = 5'b00000; w[27][123] = 5'b01111; w[27][124] = 5'b01111; w[27][125] = 5'b01111; w[27][126] = 5'b01111; w[27][127] = 5'b01111; w[27][128] = 5'b01111; w[27][129] = 5'b00000; w[27][130] = 5'b01111; w[27][131] = 5'b01111; w[27][132] = 5'b00000; w[27][133] = 5'b10000; w[27][134] = 5'b01111; w[27][135] = 5'b01111; w[27][136] = 5'b00000; w[27][137] = 5'b01111; w[27][138] = 5'b01111; w[27][139] = 5'b01111; w[27][140] = 5'b01111; w[27][141] = 5'b01111; w[27][142] = 5'b01111; w[27][143] = 5'b00000; w[27][144] = 5'b00000; w[27][145] = 5'b01111; w[27][146] = 5'b00000; w[27][147] = 5'b10000; w[27][148] = 5'b01111; w[27][149] = 5'b00000; w[27][150] = 5'b00000; w[27][151] = 5'b01111; w[27][152] = 5'b01111; w[27][153] = 5'b01111; w[27][154] = 5'b01111; w[27][155] = 5'b01111; w[27][156] = 5'b01111; w[27][157] = 5'b00000; w[27][158] = 5'b00000; w[27][159] = 5'b00000; w[27][160] = 5'b10000; w[27][161] = 5'b10000; w[27][162] = 5'b10000; w[27][163] = 5'b00000; w[27][164] = 5'b00000; w[27][165] = 5'b01111; w[27][166] = 5'b01111; w[27][167] = 5'b01111; w[27][168] = 5'b01111; w[27][169] = 5'b01111; w[27][170] = 5'b01111; w[27][171] = 5'b01111; w[27][172] = 5'b00000; w[27][173] = 5'b00000; w[27][174] = 5'b10000; w[27][175] = 5'b10000; w[27][176] = 5'b10000; w[27][177] = 5'b00000; w[27][178] = 5'b01111; w[27][179] = 5'b01111; w[27][180] = 5'b01111; w[27][181] = 5'b01111; w[27][182] = 5'b01111; w[27][183] = 5'b01111; w[27][184] = 5'b01111; w[27][185] = 5'b01111; w[27][186] = 5'b01111; w[27][187] = 5'b01111; w[27][188] = 5'b01111; w[27][189] = 5'b01111; w[27][190] = 5'b01111; w[27][191] = 5'b01111; w[27][192] = 5'b01111; w[27][193] = 5'b01111; w[27][194] = 5'b01111; w[27][195] = 5'b01111; w[27][196] = 5'b01111; w[27][197] = 5'b01111; w[27][198] = 5'b01111; w[27][199] = 5'b01111; w[27][200] = 5'b01111; w[27][201] = 5'b01111; w[27][202] = 5'b01111; w[27][203] = 5'b01111; w[27][204] = 5'b01111; w[27][205] = 5'b01111; w[27][206] = 5'b01111; w[27][207] = 5'b01111; w[27][208] = 5'b01111; w[27][209] = 5'b01111; 
w[28][0] = 5'b01111; w[28][1] = 5'b01111; w[28][2] = 5'b01111; w[28][3] = 5'b01111; w[28][4] = 5'b01111; w[28][5] = 5'b01111; w[28][6] = 5'b01111; w[28][7] = 5'b01111; w[28][8] = 5'b01111; w[28][9] = 5'b01111; w[28][10] = 5'b01111; w[28][11] = 5'b01111; w[28][12] = 5'b01111; w[28][13] = 5'b01111; w[28][14] = 5'b01111; w[28][15] = 5'b01111; w[28][16] = 5'b01111; w[28][17] = 5'b01111; w[28][18] = 5'b01111; w[28][19] = 5'b01111; w[28][20] = 5'b01111; w[28][21] = 5'b01111; w[28][22] = 5'b01111; w[28][23] = 5'b01111; w[28][24] = 5'b01111; w[28][25] = 5'b01111; w[28][26] = 5'b01111; w[28][27] = 5'b01111; w[28][28] = 5'b00000; w[28][29] = 5'b01111; w[28][30] = 5'b01111; w[28][31] = 5'b00000; w[28][32] = 5'b10000; w[28][33] = 5'b10000; w[28][34] = 5'b10000; w[28][35] = 5'b10000; w[28][36] = 5'b10000; w[28][37] = 5'b10000; w[28][38] = 5'b00000; w[28][39] = 5'b01111; w[28][40] = 5'b01111; w[28][41] = 5'b01111; w[28][42] = 5'b01111; w[28][43] = 5'b01111; w[28][44] = 5'b01111; w[28][45] = 5'b10000; w[28][46] = 5'b10000; w[28][47] = 5'b10000; w[28][48] = 5'b10000; w[28][49] = 5'b10000; w[28][50] = 5'b10000; w[28][51] = 5'b10000; w[28][52] = 5'b10000; w[28][53] = 5'b01111; w[28][54] = 5'b01111; w[28][55] = 5'b01111; w[28][56] = 5'b01111; w[28][57] = 5'b01111; w[28][58] = 5'b01111; w[28][59] = 5'b00000; w[28][60] = 5'b00000; w[28][61] = 5'b01111; w[28][62] = 5'b10000; w[28][63] = 5'b00000; w[28][64] = 5'b01111; w[28][65] = 5'b00000; w[28][66] = 5'b00000; w[28][67] = 5'b01111; w[28][68] = 5'b01111; w[28][69] = 5'b01111; w[28][70] = 5'b01111; w[28][71] = 5'b01111; w[28][72] = 5'b01111; w[28][73] = 5'b00000; w[28][74] = 5'b01111; w[28][75] = 5'b01111; w[28][76] = 5'b10000; w[28][77] = 5'b00000; w[28][78] = 5'b01111; w[28][79] = 5'b01111; w[28][80] = 5'b00000; w[28][81] = 5'b01111; w[28][82] = 5'b01111; w[28][83] = 5'b01111; w[28][84] = 5'b01111; w[28][85] = 5'b01111; w[28][86] = 5'b01111; w[28][87] = 5'b00000; w[28][88] = 5'b01111; w[28][89] = 5'b01111; w[28][90] = 5'b10000; w[28][91] = 5'b10000; w[28][92] = 5'b01111; w[28][93] = 5'b01111; w[28][94] = 5'b01111; w[28][95] = 5'b01111; w[28][96] = 5'b01111; w[28][97] = 5'b01111; w[28][98] = 5'b01111; w[28][99] = 5'b01111; w[28][100] = 5'b01111; w[28][101] = 5'b00000; w[28][102] = 5'b01111; w[28][103] = 5'b01111; w[28][104] = 5'b10000; w[28][105] = 5'b10000; w[28][106] = 5'b01111; w[28][107] = 5'b00000; w[28][108] = 5'b00000; w[28][109] = 5'b01111; w[28][110] = 5'b01111; w[28][111] = 5'b01111; w[28][112] = 5'b01111; w[28][113] = 5'b01111; w[28][114] = 5'b01111; w[28][115] = 5'b00000; w[28][116] = 5'b01111; w[28][117] = 5'b01111; w[28][118] = 5'b10000; w[28][119] = 5'b10000; w[28][120] = 5'b00000; w[28][121] = 5'b00000; w[28][122] = 5'b00000; w[28][123] = 5'b01111; w[28][124] = 5'b01111; w[28][125] = 5'b01111; w[28][126] = 5'b01111; w[28][127] = 5'b01111; w[28][128] = 5'b01111; w[28][129] = 5'b00000; w[28][130] = 5'b01111; w[28][131] = 5'b01111; w[28][132] = 5'b00000; w[28][133] = 5'b10000; w[28][134] = 5'b01111; w[28][135] = 5'b01111; w[28][136] = 5'b00000; w[28][137] = 5'b01111; w[28][138] = 5'b01111; w[28][139] = 5'b01111; w[28][140] = 5'b01111; w[28][141] = 5'b01111; w[28][142] = 5'b01111; w[28][143] = 5'b00000; w[28][144] = 5'b00000; w[28][145] = 5'b01111; w[28][146] = 5'b00000; w[28][147] = 5'b10000; w[28][148] = 5'b01111; w[28][149] = 5'b00000; w[28][150] = 5'b00000; w[28][151] = 5'b01111; w[28][152] = 5'b01111; w[28][153] = 5'b01111; w[28][154] = 5'b01111; w[28][155] = 5'b01111; w[28][156] = 5'b01111; w[28][157] = 5'b00000; w[28][158] = 5'b00000; w[28][159] = 5'b00000; w[28][160] = 5'b10000; w[28][161] = 5'b10000; w[28][162] = 5'b10000; w[28][163] = 5'b00000; w[28][164] = 5'b00000; w[28][165] = 5'b01111; w[28][166] = 5'b01111; w[28][167] = 5'b01111; w[28][168] = 5'b01111; w[28][169] = 5'b01111; w[28][170] = 5'b01111; w[28][171] = 5'b01111; w[28][172] = 5'b00000; w[28][173] = 5'b00000; w[28][174] = 5'b10000; w[28][175] = 5'b10000; w[28][176] = 5'b10000; w[28][177] = 5'b00000; w[28][178] = 5'b01111; w[28][179] = 5'b01111; w[28][180] = 5'b01111; w[28][181] = 5'b01111; w[28][182] = 5'b01111; w[28][183] = 5'b01111; w[28][184] = 5'b01111; w[28][185] = 5'b01111; w[28][186] = 5'b01111; w[28][187] = 5'b01111; w[28][188] = 5'b01111; w[28][189] = 5'b01111; w[28][190] = 5'b01111; w[28][191] = 5'b01111; w[28][192] = 5'b01111; w[28][193] = 5'b01111; w[28][194] = 5'b01111; w[28][195] = 5'b01111; w[28][196] = 5'b01111; w[28][197] = 5'b01111; w[28][198] = 5'b01111; w[28][199] = 5'b01111; w[28][200] = 5'b01111; w[28][201] = 5'b01111; w[28][202] = 5'b01111; w[28][203] = 5'b01111; w[28][204] = 5'b01111; w[28][205] = 5'b01111; w[28][206] = 5'b01111; w[28][207] = 5'b01111; w[28][208] = 5'b01111; w[28][209] = 5'b01111; 
w[29][0] = 5'b01111; w[29][1] = 5'b01111; w[29][2] = 5'b01111; w[29][3] = 5'b01111; w[29][4] = 5'b01111; w[29][5] = 5'b01111; w[29][6] = 5'b01111; w[29][7] = 5'b01111; w[29][8] = 5'b01111; w[29][9] = 5'b01111; w[29][10] = 5'b01111; w[29][11] = 5'b01111; w[29][12] = 5'b01111; w[29][13] = 5'b01111; w[29][14] = 5'b01111; w[29][15] = 5'b01111; w[29][16] = 5'b01111; w[29][17] = 5'b01111; w[29][18] = 5'b01111; w[29][19] = 5'b01111; w[29][20] = 5'b01111; w[29][21] = 5'b01111; w[29][22] = 5'b01111; w[29][23] = 5'b01111; w[29][24] = 5'b01111; w[29][25] = 5'b01111; w[29][26] = 5'b01111; w[29][27] = 5'b01111; w[29][28] = 5'b01111; w[29][29] = 5'b00000; w[29][30] = 5'b01111; w[29][31] = 5'b00000; w[29][32] = 5'b10000; w[29][33] = 5'b10000; w[29][34] = 5'b10000; w[29][35] = 5'b10000; w[29][36] = 5'b10000; w[29][37] = 5'b10000; w[29][38] = 5'b00000; w[29][39] = 5'b01111; w[29][40] = 5'b01111; w[29][41] = 5'b01111; w[29][42] = 5'b01111; w[29][43] = 5'b01111; w[29][44] = 5'b01111; w[29][45] = 5'b10000; w[29][46] = 5'b10000; w[29][47] = 5'b10000; w[29][48] = 5'b10000; w[29][49] = 5'b10000; w[29][50] = 5'b10000; w[29][51] = 5'b10000; w[29][52] = 5'b10000; w[29][53] = 5'b01111; w[29][54] = 5'b01111; w[29][55] = 5'b01111; w[29][56] = 5'b01111; w[29][57] = 5'b01111; w[29][58] = 5'b01111; w[29][59] = 5'b00000; w[29][60] = 5'b00000; w[29][61] = 5'b01111; w[29][62] = 5'b10000; w[29][63] = 5'b00000; w[29][64] = 5'b01111; w[29][65] = 5'b00000; w[29][66] = 5'b00000; w[29][67] = 5'b01111; w[29][68] = 5'b01111; w[29][69] = 5'b01111; w[29][70] = 5'b01111; w[29][71] = 5'b01111; w[29][72] = 5'b01111; w[29][73] = 5'b00000; w[29][74] = 5'b01111; w[29][75] = 5'b01111; w[29][76] = 5'b10000; w[29][77] = 5'b00000; w[29][78] = 5'b01111; w[29][79] = 5'b01111; w[29][80] = 5'b00000; w[29][81] = 5'b01111; w[29][82] = 5'b01111; w[29][83] = 5'b01111; w[29][84] = 5'b01111; w[29][85] = 5'b01111; w[29][86] = 5'b01111; w[29][87] = 5'b00000; w[29][88] = 5'b01111; w[29][89] = 5'b01111; w[29][90] = 5'b10000; w[29][91] = 5'b10000; w[29][92] = 5'b01111; w[29][93] = 5'b01111; w[29][94] = 5'b01111; w[29][95] = 5'b01111; w[29][96] = 5'b01111; w[29][97] = 5'b01111; w[29][98] = 5'b01111; w[29][99] = 5'b01111; w[29][100] = 5'b01111; w[29][101] = 5'b00000; w[29][102] = 5'b01111; w[29][103] = 5'b01111; w[29][104] = 5'b10000; w[29][105] = 5'b10000; w[29][106] = 5'b01111; w[29][107] = 5'b00000; w[29][108] = 5'b00000; w[29][109] = 5'b01111; w[29][110] = 5'b01111; w[29][111] = 5'b01111; w[29][112] = 5'b01111; w[29][113] = 5'b01111; w[29][114] = 5'b01111; w[29][115] = 5'b00000; w[29][116] = 5'b01111; w[29][117] = 5'b01111; w[29][118] = 5'b10000; w[29][119] = 5'b10000; w[29][120] = 5'b00000; w[29][121] = 5'b00000; w[29][122] = 5'b00000; w[29][123] = 5'b01111; w[29][124] = 5'b01111; w[29][125] = 5'b01111; w[29][126] = 5'b01111; w[29][127] = 5'b01111; w[29][128] = 5'b01111; w[29][129] = 5'b00000; w[29][130] = 5'b01111; w[29][131] = 5'b01111; w[29][132] = 5'b00000; w[29][133] = 5'b10000; w[29][134] = 5'b01111; w[29][135] = 5'b01111; w[29][136] = 5'b00000; w[29][137] = 5'b01111; w[29][138] = 5'b01111; w[29][139] = 5'b01111; w[29][140] = 5'b01111; w[29][141] = 5'b01111; w[29][142] = 5'b01111; w[29][143] = 5'b00000; w[29][144] = 5'b00000; w[29][145] = 5'b01111; w[29][146] = 5'b00000; w[29][147] = 5'b10000; w[29][148] = 5'b01111; w[29][149] = 5'b00000; w[29][150] = 5'b00000; w[29][151] = 5'b01111; w[29][152] = 5'b01111; w[29][153] = 5'b01111; w[29][154] = 5'b01111; w[29][155] = 5'b01111; w[29][156] = 5'b01111; w[29][157] = 5'b00000; w[29][158] = 5'b00000; w[29][159] = 5'b00000; w[29][160] = 5'b10000; w[29][161] = 5'b10000; w[29][162] = 5'b10000; w[29][163] = 5'b00000; w[29][164] = 5'b00000; w[29][165] = 5'b01111; w[29][166] = 5'b01111; w[29][167] = 5'b01111; w[29][168] = 5'b01111; w[29][169] = 5'b01111; w[29][170] = 5'b01111; w[29][171] = 5'b01111; w[29][172] = 5'b00000; w[29][173] = 5'b00000; w[29][174] = 5'b10000; w[29][175] = 5'b10000; w[29][176] = 5'b10000; w[29][177] = 5'b00000; w[29][178] = 5'b01111; w[29][179] = 5'b01111; w[29][180] = 5'b01111; w[29][181] = 5'b01111; w[29][182] = 5'b01111; w[29][183] = 5'b01111; w[29][184] = 5'b01111; w[29][185] = 5'b01111; w[29][186] = 5'b01111; w[29][187] = 5'b01111; w[29][188] = 5'b01111; w[29][189] = 5'b01111; w[29][190] = 5'b01111; w[29][191] = 5'b01111; w[29][192] = 5'b01111; w[29][193] = 5'b01111; w[29][194] = 5'b01111; w[29][195] = 5'b01111; w[29][196] = 5'b01111; w[29][197] = 5'b01111; w[29][198] = 5'b01111; w[29][199] = 5'b01111; w[29][200] = 5'b01111; w[29][201] = 5'b01111; w[29][202] = 5'b01111; w[29][203] = 5'b01111; w[29][204] = 5'b01111; w[29][205] = 5'b01111; w[29][206] = 5'b01111; w[29][207] = 5'b01111; w[29][208] = 5'b01111; w[29][209] = 5'b01111; 
w[30][0] = 5'b01111; w[30][1] = 5'b01111; w[30][2] = 5'b01111; w[30][3] = 5'b01111; w[30][4] = 5'b01111; w[30][5] = 5'b01111; w[30][6] = 5'b01111; w[30][7] = 5'b01111; w[30][8] = 5'b01111; w[30][9] = 5'b01111; w[30][10] = 5'b01111; w[30][11] = 5'b01111; w[30][12] = 5'b01111; w[30][13] = 5'b01111; w[30][14] = 5'b01111; w[30][15] = 5'b01111; w[30][16] = 5'b01111; w[30][17] = 5'b01111; w[30][18] = 5'b01111; w[30][19] = 5'b01111; w[30][20] = 5'b01111; w[30][21] = 5'b01111; w[30][22] = 5'b01111; w[30][23] = 5'b01111; w[30][24] = 5'b01111; w[30][25] = 5'b01111; w[30][26] = 5'b01111; w[30][27] = 5'b01111; w[30][28] = 5'b01111; w[30][29] = 5'b01111; w[30][30] = 5'b00000; w[30][31] = 5'b01111; w[30][32] = 5'b00000; w[30][33] = 5'b10000; w[30][34] = 5'b00000; w[30][35] = 5'b00000; w[30][36] = 5'b00000; w[30][37] = 5'b00000; w[30][38] = 5'b01111; w[30][39] = 5'b01111; w[30][40] = 5'b01111; w[30][41] = 5'b01111; w[30][42] = 5'b01111; w[30][43] = 5'b01111; w[30][44] = 5'b01111; w[30][45] = 5'b00000; w[30][46] = 5'b00000; w[30][47] = 5'b10000; w[30][48] = 5'b00000; w[30][49] = 5'b00000; w[30][50] = 5'b00000; w[30][51] = 5'b00000; w[30][52] = 5'b00000; w[30][53] = 5'b01111; w[30][54] = 5'b01111; w[30][55] = 5'b01111; w[30][56] = 5'b01111; w[30][57] = 5'b01111; w[30][58] = 5'b00000; w[30][59] = 5'b10000; w[30][60] = 5'b10000; w[30][61] = 5'b00000; w[30][62] = 5'b00000; w[30][63] = 5'b01111; w[30][64] = 5'b01111; w[30][65] = 5'b10000; w[30][66] = 5'b10000; w[30][67] = 5'b00000; w[30][68] = 5'b01111; w[30][69] = 5'b01111; w[30][70] = 5'b01111; w[30][71] = 5'b01111; w[30][72] = 5'b00000; w[30][73] = 5'b10000; w[30][74] = 5'b00000; w[30][75] = 5'b00000; w[30][76] = 5'b00000; w[30][77] = 5'b01111; w[30][78] = 5'b01111; w[30][79] = 5'b00000; w[30][80] = 5'b10000; w[30][81] = 5'b00000; w[30][82] = 5'b01111; w[30][83] = 5'b01111; w[30][84] = 5'b01111; w[30][85] = 5'b01111; w[30][86] = 5'b00000; w[30][87] = 5'b10000; w[30][88] = 5'b00000; w[30][89] = 5'b00000; w[30][90] = 5'b00000; w[30][91] = 5'b00000; w[30][92] = 5'b01111; w[30][93] = 5'b00000; w[30][94] = 5'b00000; w[30][95] = 5'b01111; w[30][96] = 5'b01111; w[30][97] = 5'b01111; w[30][98] = 5'b01111; w[30][99] = 5'b01111; w[30][100] = 5'b00000; w[30][101] = 5'b10000; w[30][102] = 5'b00000; w[30][103] = 5'b01111; w[30][104] = 5'b00000; w[30][105] = 5'b00000; w[30][106] = 5'b00000; w[30][107] = 5'b10000; w[30][108] = 5'b10000; w[30][109] = 5'b00000; w[30][110] = 5'b01111; w[30][111] = 5'b01111; w[30][112] = 5'b01111; w[30][113] = 5'b01111; w[30][114] = 5'b00000; w[30][115] = 5'b10000; w[30][116] = 5'b00000; w[30][117] = 5'b01111; w[30][118] = 5'b00000; w[30][119] = 5'b00000; w[30][120] = 5'b10000; w[30][121] = 5'b10000; w[30][122] = 5'b10000; w[30][123] = 5'b00000; w[30][124] = 5'b01111; w[30][125] = 5'b01111; w[30][126] = 5'b01111; w[30][127] = 5'b01111; w[30][128] = 5'b00000; w[30][129] = 5'b10000; w[30][130] = 5'b00000; w[30][131] = 5'b01111; w[30][132] = 5'b01111; w[30][133] = 5'b00000; w[30][134] = 5'b00000; w[30][135] = 5'b00000; w[30][136] = 5'b10000; w[30][137] = 5'b00000; w[30][138] = 5'b01111; w[30][139] = 5'b01111; w[30][140] = 5'b01111; w[30][141] = 5'b01111; w[30][142] = 5'b00000; w[30][143] = 5'b10000; w[30][144] = 5'b10000; w[30][145] = 5'b01111; w[30][146] = 5'b01111; w[30][147] = 5'b00000; w[30][148] = 5'b00000; w[30][149] = 5'b10000; w[30][150] = 5'b10000; w[30][151] = 5'b00000; w[30][152] = 5'b01111; w[30][153] = 5'b01111; w[30][154] = 5'b01111; w[30][155] = 5'b01111; w[30][156] = 5'b01111; w[30][157] = 5'b10000; w[30][158] = 5'b10000; w[30][159] = 5'b10000; w[30][160] = 5'b00000; w[30][161] = 5'b00000; w[30][162] = 5'b10000; w[30][163] = 5'b10000; w[30][164] = 5'b10000; w[30][165] = 5'b01111; w[30][166] = 5'b01111; w[30][167] = 5'b01111; w[30][168] = 5'b01111; w[30][169] = 5'b01111; w[30][170] = 5'b01111; w[30][171] = 5'b00000; w[30][172] = 5'b10000; w[30][173] = 5'b10000; w[30][174] = 5'b00000; w[30][175] = 5'b00000; w[30][176] = 5'b10000; w[30][177] = 5'b10000; w[30][178] = 5'b00000; w[30][179] = 5'b01111; w[30][180] = 5'b01111; w[30][181] = 5'b01111; w[30][182] = 5'b01111; w[30][183] = 5'b01111; w[30][184] = 5'b01111; w[30][185] = 5'b01111; w[30][186] = 5'b01111; w[30][187] = 5'b01111; w[30][188] = 5'b01111; w[30][189] = 5'b01111; w[30][190] = 5'b01111; w[30][191] = 5'b01111; w[30][192] = 5'b01111; w[30][193] = 5'b01111; w[30][194] = 5'b01111; w[30][195] = 5'b01111; w[30][196] = 5'b01111; w[30][197] = 5'b01111; w[30][198] = 5'b01111; w[30][199] = 5'b01111; w[30][200] = 5'b01111; w[30][201] = 5'b01111; w[30][202] = 5'b01111; w[30][203] = 5'b01111; w[30][204] = 5'b01111; w[30][205] = 5'b01111; w[30][206] = 5'b01111; w[30][207] = 5'b01111; w[30][208] = 5'b01111; w[30][209] = 5'b01111; 
w[31][0] = 5'b00000; w[31][1] = 5'b00000; w[31][2] = 5'b00000; w[31][3] = 5'b00000; w[31][4] = 5'b00000; w[31][5] = 5'b00000; w[31][6] = 5'b00000; w[31][7] = 5'b00000; w[31][8] = 5'b00000; w[31][9] = 5'b00000; w[31][10] = 5'b00000; w[31][11] = 5'b00000; w[31][12] = 5'b00000; w[31][13] = 5'b00000; w[31][14] = 5'b00000; w[31][15] = 5'b00000; w[31][16] = 5'b00000; w[31][17] = 5'b00000; w[31][18] = 5'b00000; w[31][19] = 5'b00000; w[31][20] = 5'b00000; w[31][21] = 5'b00000; w[31][22] = 5'b00000; w[31][23] = 5'b00000; w[31][24] = 5'b00000; w[31][25] = 5'b00000; w[31][26] = 5'b00000; w[31][27] = 5'b00000; w[31][28] = 5'b00000; w[31][29] = 5'b00000; w[31][30] = 5'b01111; w[31][31] = 5'b00000; w[31][32] = 5'b01111; w[31][33] = 5'b00000; w[31][34] = 5'b10000; w[31][35] = 5'b10000; w[31][36] = 5'b10000; w[31][37] = 5'b01111; w[31][38] = 5'b01111; w[31][39] = 5'b01111; w[31][40] = 5'b00000; w[31][41] = 5'b00000; w[31][42] = 5'b00000; w[31][43] = 5'b00000; w[31][44] = 5'b01111; w[31][45] = 5'b01111; w[31][46] = 5'b01111; w[31][47] = 5'b00000; w[31][48] = 5'b10000; w[31][49] = 5'b10000; w[31][50] = 5'b10000; w[31][51] = 5'b01111; w[31][52] = 5'b01111; w[31][53] = 5'b01111; w[31][54] = 5'b00000; w[31][55] = 5'b00000; w[31][56] = 5'b00000; w[31][57] = 5'b00000; w[31][58] = 5'b10000; w[31][59] = 5'b00000; w[31][60] = 5'b00000; w[31][61] = 5'b01111; w[31][62] = 5'b01111; w[31][63] = 5'b00000; w[31][64] = 5'b00000; w[31][65] = 5'b00000; w[31][66] = 5'b00000; w[31][67] = 5'b10000; w[31][68] = 5'b00000; w[31][69] = 5'b00000; w[31][70] = 5'b00000; w[31][71] = 5'b00000; w[31][72] = 5'b10000; w[31][73] = 5'b00000; w[31][74] = 5'b01111; w[31][75] = 5'b01111; w[31][76] = 5'b01111; w[31][77] = 5'b00000; w[31][78] = 5'b00000; w[31][79] = 5'b01111; w[31][80] = 5'b00000; w[31][81] = 5'b10000; w[31][82] = 5'b00000; w[31][83] = 5'b00000; w[31][84] = 5'b00000; w[31][85] = 5'b00000; w[31][86] = 5'b10000; w[31][87] = 5'b00000; w[31][88] = 5'b01111; w[31][89] = 5'b01111; w[31][90] = 5'b01111; w[31][91] = 5'b01111; w[31][92] = 5'b00000; w[31][93] = 5'b01111; w[31][94] = 5'b01111; w[31][95] = 5'b00000; w[31][96] = 5'b00000; w[31][97] = 5'b00000; w[31][98] = 5'b00000; w[31][99] = 5'b00000; w[31][100] = 5'b10000; w[31][101] = 5'b00000; w[31][102] = 5'b01111; w[31][103] = 5'b00000; w[31][104] = 5'b01111; w[31][105] = 5'b01111; w[31][106] = 5'b10000; w[31][107] = 5'b00000; w[31][108] = 5'b00000; w[31][109] = 5'b10000; w[31][110] = 5'b00000; w[31][111] = 5'b00000; w[31][112] = 5'b00000; w[31][113] = 5'b00000; w[31][114] = 5'b10000; w[31][115] = 5'b00000; w[31][116] = 5'b01111; w[31][117] = 5'b00000; w[31][118] = 5'b01111; w[31][119] = 5'b01111; w[31][120] = 5'b00000; w[31][121] = 5'b00000; w[31][122] = 5'b00000; w[31][123] = 5'b10000; w[31][124] = 5'b00000; w[31][125] = 5'b00000; w[31][126] = 5'b00000; w[31][127] = 5'b00000; w[31][128] = 5'b10000; w[31][129] = 5'b00000; w[31][130] = 5'b01111; w[31][131] = 5'b00000; w[31][132] = 5'b00000; w[31][133] = 5'b01111; w[31][134] = 5'b01111; w[31][135] = 5'b01111; w[31][136] = 5'b00000; w[31][137] = 5'b10000; w[31][138] = 5'b00000; w[31][139] = 5'b00000; w[31][140] = 5'b00000; w[31][141] = 5'b00000; w[31][142] = 5'b10000; w[31][143] = 5'b00000; w[31][144] = 5'b00000; w[31][145] = 5'b00000; w[31][146] = 5'b00000; w[31][147] = 5'b01111; w[31][148] = 5'b01111; w[31][149] = 5'b00000; w[31][150] = 5'b00000; w[31][151] = 5'b10000; w[31][152] = 5'b00000; w[31][153] = 5'b00000; w[31][154] = 5'b00000; w[31][155] = 5'b00000; w[31][156] = 5'b00000; w[31][157] = 5'b00000; w[31][158] = 5'b00000; w[31][159] = 5'b10000; w[31][160] = 5'b10000; w[31][161] = 5'b10000; w[31][162] = 5'b10000; w[31][163] = 5'b00000; w[31][164] = 5'b00000; w[31][165] = 5'b00000; w[31][166] = 5'b00000; w[31][167] = 5'b00000; w[31][168] = 5'b00000; w[31][169] = 5'b00000; w[31][170] = 5'b00000; w[31][171] = 5'b01111; w[31][172] = 5'b00000; w[31][173] = 5'b10000; w[31][174] = 5'b10000; w[31][175] = 5'b10000; w[31][176] = 5'b10000; w[31][177] = 5'b00000; w[31][178] = 5'b01111; w[31][179] = 5'b00000; w[31][180] = 5'b00000; w[31][181] = 5'b00000; w[31][182] = 5'b00000; w[31][183] = 5'b00000; w[31][184] = 5'b00000; w[31][185] = 5'b00000; w[31][186] = 5'b00000; w[31][187] = 5'b00000; w[31][188] = 5'b00000; w[31][189] = 5'b00000; w[31][190] = 5'b00000; w[31][191] = 5'b00000; w[31][192] = 5'b00000; w[31][193] = 5'b00000; w[31][194] = 5'b00000; w[31][195] = 5'b00000; w[31][196] = 5'b00000; w[31][197] = 5'b00000; w[31][198] = 5'b00000; w[31][199] = 5'b00000; w[31][200] = 5'b00000; w[31][201] = 5'b00000; w[31][202] = 5'b00000; w[31][203] = 5'b00000; w[31][204] = 5'b00000; w[31][205] = 5'b00000; w[31][206] = 5'b00000; w[31][207] = 5'b00000; w[31][208] = 5'b00000; w[31][209] = 5'b00000; 
w[32][0] = 5'b10000; w[32][1] = 5'b10000; w[32][2] = 5'b10000; w[32][3] = 5'b10000; w[32][4] = 5'b10000; w[32][5] = 5'b10000; w[32][6] = 5'b10000; w[32][7] = 5'b10000; w[32][8] = 5'b10000; w[32][9] = 5'b10000; w[32][10] = 5'b10000; w[32][11] = 5'b10000; w[32][12] = 5'b10000; w[32][13] = 5'b10000; w[32][14] = 5'b10000; w[32][15] = 5'b10000; w[32][16] = 5'b10000; w[32][17] = 5'b10000; w[32][18] = 5'b10000; w[32][19] = 5'b10000; w[32][20] = 5'b10000; w[32][21] = 5'b10000; w[32][22] = 5'b10000; w[32][23] = 5'b10000; w[32][24] = 5'b10000; w[32][25] = 5'b10000; w[32][26] = 5'b10000; w[32][27] = 5'b10000; w[32][28] = 5'b10000; w[32][29] = 5'b10000; w[32][30] = 5'b00000; w[32][31] = 5'b01111; w[32][32] = 5'b00000; w[32][33] = 5'b01111; w[32][34] = 5'b00000; w[32][35] = 5'b00000; w[32][36] = 5'b00000; w[32][37] = 5'b01111; w[32][38] = 5'b01111; w[32][39] = 5'b00000; w[32][40] = 5'b10000; w[32][41] = 5'b10000; w[32][42] = 5'b10000; w[32][43] = 5'b10000; w[32][44] = 5'b00000; w[32][45] = 5'b01111; w[32][46] = 5'b01111; w[32][47] = 5'b01111; w[32][48] = 5'b00000; w[32][49] = 5'b00000; w[32][50] = 5'b00000; w[32][51] = 5'b01111; w[32][52] = 5'b01111; w[32][53] = 5'b00000; w[32][54] = 5'b10000; w[32][55] = 5'b10000; w[32][56] = 5'b10000; w[32][57] = 5'b10000; w[32][58] = 5'b00000; w[32][59] = 5'b01111; w[32][60] = 5'b01111; w[32][61] = 5'b00000; w[32][62] = 5'b00000; w[32][63] = 5'b10000; w[32][64] = 5'b10000; w[32][65] = 5'b01111; w[32][66] = 5'b01111; w[32][67] = 5'b00000; w[32][68] = 5'b10000; w[32][69] = 5'b10000; w[32][70] = 5'b10000; w[32][71] = 5'b10000; w[32][72] = 5'b00000; w[32][73] = 5'b01111; w[32][74] = 5'b00000; w[32][75] = 5'b00000; w[32][76] = 5'b00000; w[32][77] = 5'b10000; w[32][78] = 5'b10000; w[32][79] = 5'b00000; w[32][80] = 5'b01111; w[32][81] = 5'b00000; w[32][82] = 5'b10000; w[32][83] = 5'b10000; w[32][84] = 5'b10000; w[32][85] = 5'b10000; w[32][86] = 5'b00000; w[32][87] = 5'b01111; w[32][88] = 5'b00000; w[32][89] = 5'b00000; w[32][90] = 5'b00000; w[32][91] = 5'b00000; w[32][92] = 5'b10000; w[32][93] = 5'b00000; w[32][94] = 5'b00000; w[32][95] = 5'b10000; w[32][96] = 5'b10000; w[32][97] = 5'b10000; w[32][98] = 5'b10000; w[32][99] = 5'b10000; w[32][100] = 5'b00000; w[32][101] = 5'b01111; w[32][102] = 5'b00000; w[32][103] = 5'b10000; w[32][104] = 5'b00000; w[32][105] = 5'b00000; w[32][106] = 5'b00000; w[32][107] = 5'b01111; w[32][108] = 5'b01111; w[32][109] = 5'b00000; w[32][110] = 5'b10000; w[32][111] = 5'b10000; w[32][112] = 5'b10000; w[32][113] = 5'b10000; w[32][114] = 5'b00000; w[32][115] = 5'b01111; w[32][116] = 5'b00000; w[32][117] = 5'b10000; w[32][118] = 5'b00000; w[32][119] = 5'b00000; w[32][120] = 5'b01111; w[32][121] = 5'b01111; w[32][122] = 5'b01111; w[32][123] = 5'b00000; w[32][124] = 5'b10000; w[32][125] = 5'b10000; w[32][126] = 5'b10000; w[32][127] = 5'b10000; w[32][128] = 5'b00000; w[32][129] = 5'b01111; w[32][130] = 5'b00000; w[32][131] = 5'b10000; w[32][132] = 5'b10000; w[32][133] = 5'b00000; w[32][134] = 5'b00000; w[32][135] = 5'b00000; w[32][136] = 5'b01111; w[32][137] = 5'b00000; w[32][138] = 5'b10000; w[32][139] = 5'b10000; w[32][140] = 5'b10000; w[32][141] = 5'b10000; w[32][142] = 5'b00000; w[32][143] = 5'b01111; w[32][144] = 5'b01111; w[32][145] = 5'b10000; w[32][146] = 5'b10000; w[32][147] = 5'b00000; w[32][148] = 5'b00000; w[32][149] = 5'b01111; w[32][150] = 5'b01111; w[32][151] = 5'b00000; w[32][152] = 5'b10000; w[32][153] = 5'b10000; w[32][154] = 5'b10000; w[32][155] = 5'b10000; w[32][156] = 5'b10000; w[32][157] = 5'b01111; w[32][158] = 5'b01111; w[32][159] = 5'b10000; w[32][160] = 5'b00000; w[32][161] = 5'b00000; w[32][162] = 5'b00000; w[32][163] = 5'b01111; w[32][164] = 5'b01111; w[32][165] = 5'b10000; w[32][166] = 5'b10000; w[32][167] = 5'b10000; w[32][168] = 5'b10000; w[32][169] = 5'b10000; w[32][170] = 5'b10000; w[32][171] = 5'b00000; w[32][172] = 5'b01111; w[32][173] = 5'b10000; w[32][174] = 5'b00000; w[32][175] = 5'b00000; w[32][176] = 5'b00000; w[32][177] = 5'b01111; w[32][178] = 5'b00000; w[32][179] = 5'b10000; w[32][180] = 5'b10000; w[32][181] = 5'b10000; w[32][182] = 5'b10000; w[32][183] = 5'b10000; w[32][184] = 5'b10000; w[32][185] = 5'b10000; w[32][186] = 5'b10000; w[32][187] = 5'b10000; w[32][188] = 5'b10000; w[32][189] = 5'b10000; w[32][190] = 5'b10000; w[32][191] = 5'b10000; w[32][192] = 5'b10000; w[32][193] = 5'b10000; w[32][194] = 5'b10000; w[32][195] = 5'b10000; w[32][196] = 5'b10000; w[32][197] = 5'b10000; w[32][198] = 5'b10000; w[32][199] = 5'b10000; w[32][200] = 5'b10000; w[32][201] = 5'b10000; w[32][202] = 5'b10000; w[32][203] = 5'b10000; w[32][204] = 5'b10000; w[32][205] = 5'b10000; w[32][206] = 5'b10000; w[32][207] = 5'b10000; w[32][208] = 5'b10000; w[32][209] = 5'b10000; 
w[33][0] = 5'b10000; w[33][1] = 5'b10000; w[33][2] = 5'b10000; w[33][3] = 5'b10000; w[33][4] = 5'b10000; w[33][5] = 5'b10000; w[33][6] = 5'b10000; w[33][7] = 5'b10000; w[33][8] = 5'b10000; w[33][9] = 5'b10000; w[33][10] = 5'b10000; w[33][11] = 5'b10000; w[33][12] = 5'b10000; w[33][13] = 5'b10000; w[33][14] = 5'b10000; w[33][15] = 5'b10000; w[33][16] = 5'b10000; w[33][17] = 5'b10000; w[33][18] = 5'b10000; w[33][19] = 5'b10000; w[33][20] = 5'b10000; w[33][21] = 5'b10000; w[33][22] = 5'b10000; w[33][23] = 5'b10000; w[33][24] = 5'b10000; w[33][25] = 5'b10000; w[33][26] = 5'b10000; w[33][27] = 5'b10000; w[33][28] = 5'b10000; w[33][29] = 5'b10000; w[33][30] = 5'b10000; w[33][31] = 5'b00000; w[33][32] = 5'b01111; w[33][33] = 5'b00000; w[33][34] = 5'b01111; w[33][35] = 5'b01111; w[33][36] = 5'b01111; w[33][37] = 5'b01111; w[33][38] = 5'b00000; w[33][39] = 5'b10000; w[33][40] = 5'b10000; w[33][41] = 5'b10000; w[33][42] = 5'b10000; w[33][43] = 5'b10000; w[33][44] = 5'b10000; w[33][45] = 5'b01111; w[33][46] = 5'b01111; w[33][47] = 5'b01111; w[33][48] = 5'b01111; w[33][49] = 5'b01111; w[33][50] = 5'b01111; w[33][51] = 5'b01111; w[33][52] = 5'b01111; w[33][53] = 5'b10000; w[33][54] = 5'b10000; w[33][55] = 5'b10000; w[33][56] = 5'b10000; w[33][57] = 5'b10000; w[33][58] = 5'b10000; w[33][59] = 5'b00000; w[33][60] = 5'b00000; w[33][61] = 5'b10000; w[33][62] = 5'b01111; w[33][63] = 5'b00000; w[33][64] = 5'b10000; w[33][65] = 5'b00000; w[33][66] = 5'b00000; w[33][67] = 5'b10000; w[33][68] = 5'b10000; w[33][69] = 5'b10000; w[33][70] = 5'b10000; w[33][71] = 5'b10000; w[33][72] = 5'b10000; w[33][73] = 5'b00000; w[33][74] = 5'b10000; w[33][75] = 5'b10000; w[33][76] = 5'b01111; w[33][77] = 5'b00000; w[33][78] = 5'b10000; w[33][79] = 5'b10000; w[33][80] = 5'b00000; w[33][81] = 5'b10000; w[33][82] = 5'b10000; w[33][83] = 5'b10000; w[33][84] = 5'b10000; w[33][85] = 5'b10000; w[33][86] = 5'b10000; w[33][87] = 5'b00000; w[33][88] = 5'b10000; w[33][89] = 5'b10000; w[33][90] = 5'b01111; w[33][91] = 5'b01111; w[33][92] = 5'b10000; w[33][93] = 5'b10000; w[33][94] = 5'b10000; w[33][95] = 5'b10000; w[33][96] = 5'b10000; w[33][97] = 5'b10000; w[33][98] = 5'b10000; w[33][99] = 5'b10000; w[33][100] = 5'b10000; w[33][101] = 5'b00000; w[33][102] = 5'b10000; w[33][103] = 5'b10000; w[33][104] = 5'b01111; w[33][105] = 5'b01111; w[33][106] = 5'b10000; w[33][107] = 5'b00000; w[33][108] = 5'b00000; w[33][109] = 5'b10000; w[33][110] = 5'b10000; w[33][111] = 5'b10000; w[33][112] = 5'b10000; w[33][113] = 5'b10000; w[33][114] = 5'b10000; w[33][115] = 5'b00000; w[33][116] = 5'b10000; w[33][117] = 5'b10000; w[33][118] = 5'b01111; w[33][119] = 5'b01111; w[33][120] = 5'b00000; w[33][121] = 5'b00000; w[33][122] = 5'b00000; w[33][123] = 5'b10000; w[33][124] = 5'b10000; w[33][125] = 5'b10000; w[33][126] = 5'b10000; w[33][127] = 5'b10000; w[33][128] = 5'b10000; w[33][129] = 5'b00000; w[33][130] = 5'b10000; w[33][131] = 5'b10000; w[33][132] = 5'b00000; w[33][133] = 5'b01111; w[33][134] = 5'b10000; w[33][135] = 5'b10000; w[33][136] = 5'b00000; w[33][137] = 5'b10000; w[33][138] = 5'b10000; w[33][139] = 5'b10000; w[33][140] = 5'b10000; w[33][141] = 5'b10000; w[33][142] = 5'b10000; w[33][143] = 5'b00000; w[33][144] = 5'b00000; w[33][145] = 5'b10000; w[33][146] = 5'b00000; w[33][147] = 5'b01111; w[33][148] = 5'b10000; w[33][149] = 5'b00000; w[33][150] = 5'b00000; w[33][151] = 5'b10000; w[33][152] = 5'b10000; w[33][153] = 5'b10000; w[33][154] = 5'b10000; w[33][155] = 5'b10000; w[33][156] = 5'b10000; w[33][157] = 5'b00000; w[33][158] = 5'b00000; w[33][159] = 5'b00000; w[33][160] = 5'b01111; w[33][161] = 5'b01111; w[33][162] = 5'b01111; w[33][163] = 5'b00000; w[33][164] = 5'b00000; w[33][165] = 5'b10000; w[33][166] = 5'b10000; w[33][167] = 5'b10000; w[33][168] = 5'b10000; w[33][169] = 5'b10000; w[33][170] = 5'b10000; w[33][171] = 5'b10000; w[33][172] = 5'b00000; w[33][173] = 5'b00000; w[33][174] = 5'b01111; w[33][175] = 5'b01111; w[33][176] = 5'b01111; w[33][177] = 5'b00000; w[33][178] = 5'b10000; w[33][179] = 5'b10000; w[33][180] = 5'b10000; w[33][181] = 5'b10000; w[33][182] = 5'b10000; w[33][183] = 5'b10000; w[33][184] = 5'b10000; w[33][185] = 5'b10000; w[33][186] = 5'b10000; w[33][187] = 5'b10000; w[33][188] = 5'b10000; w[33][189] = 5'b10000; w[33][190] = 5'b10000; w[33][191] = 5'b10000; w[33][192] = 5'b10000; w[33][193] = 5'b10000; w[33][194] = 5'b10000; w[33][195] = 5'b10000; w[33][196] = 5'b10000; w[33][197] = 5'b10000; w[33][198] = 5'b10000; w[33][199] = 5'b10000; w[33][200] = 5'b10000; w[33][201] = 5'b10000; w[33][202] = 5'b10000; w[33][203] = 5'b10000; w[33][204] = 5'b10000; w[33][205] = 5'b10000; w[33][206] = 5'b10000; w[33][207] = 5'b10000; w[33][208] = 5'b10000; w[33][209] = 5'b10000; 
w[34][0] = 5'b10000; w[34][1] = 5'b10000; w[34][2] = 5'b10000; w[34][3] = 5'b10000; w[34][4] = 5'b10000; w[34][5] = 5'b10000; w[34][6] = 5'b10000; w[34][7] = 5'b10000; w[34][8] = 5'b10000; w[34][9] = 5'b10000; w[34][10] = 5'b10000; w[34][11] = 5'b10000; w[34][12] = 5'b10000; w[34][13] = 5'b10000; w[34][14] = 5'b10000; w[34][15] = 5'b10000; w[34][16] = 5'b10000; w[34][17] = 5'b10000; w[34][18] = 5'b10000; w[34][19] = 5'b10000; w[34][20] = 5'b10000; w[34][21] = 5'b10000; w[34][22] = 5'b10000; w[34][23] = 5'b10000; w[34][24] = 5'b10000; w[34][25] = 5'b10000; w[34][26] = 5'b10000; w[34][27] = 5'b10000; w[34][28] = 5'b10000; w[34][29] = 5'b10000; w[34][30] = 5'b00000; w[34][31] = 5'b10000; w[34][32] = 5'b00000; w[34][33] = 5'b01111; w[34][34] = 5'b00000; w[34][35] = 5'b01111; w[34][36] = 5'b01111; w[34][37] = 5'b00000; w[34][38] = 5'b10000; w[34][39] = 5'b00000; w[34][40] = 5'b10000; w[34][41] = 5'b10000; w[34][42] = 5'b10000; w[34][43] = 5'b10000; w[34][44] = 5'b00000; w[34][45] = 5'b00000; w[34][46] = 5'b00000; w[34][47] = 5'b01111; w[34][48] = 5'b01111; w[34][49] = 5'b01111; w[34][50] = 5'b01111; w[34][51] = 5'b00000; w[34][52] = 5'b00000; w[34][53] = 5'b00000; w[34][54] = 5'b10000; w[34][55] = 5'b10000; w[34][56] = 5'b10000; w[34][57] = 5'b10000; w[34][58] = 5'b00000; w[34][59] = 5'b10000; w[34][60] = 5'b10000; w[34][61] = 5'b10000; w[34][62] = 5'b00000; w[34][63] = 5'b01111; w[34][64] = 5'b10000; w[34][65] = 5'b10000; w[34][66] = 5'b10000; w[34][67] = 5'b00000; w[34][68] = 5'b10000; w[34][69] = 5'b10000; w[34][70] = 5'b10000; w[34][71] = 5'b10000; w[34][72] = 5'b00000; w[34][73] = 5'b10000; w[34][74] = 5'b10000; w[34][75] = 5'b10000; w[34][76] = 5'b00000; w[34][77] = 5'b01111; w[34][78] = 5'b10000; w[34][79] = 5'b10000; w[34][80] = 5'b10000; w[34][81] = 5'b00000; w[34][82] = 5'b10000; w[34][83] = 5'b10000; w[34][84] = 5'b10000; w[34][85] = 5'b10000; w[34][86] = 5'b00000; w[34][87] = 5'b10000; w[34][88] = 5'b10000; w[34][89] = 5'b10000; w[34][90] = 5'b00000; w[34][91] = 5'b00000; w[34][92] = 5'b10000; w[34][93] = 5'b10000; w[34][94] = 5'b10000; w[34][95] = 5'b10000; w[34][96] = 5'b10000; w[34][97] = 5'b10000; w[34][98] = 5'b10000; w[34][99] = 5'b10000; w[34][100] = 5'b00000; w[34][101] = 5'b10000; w[34][102] = 5'b10000; w[34][103] = 5'b10000; w[34][104] = 5'b00000; w[34][105] = 5'b00000; w[34][106] = 5'b00000; w[34][107] = 5'b10000; w[34][108] = 5'b10000; w[34][109] = 5'b00000; w[34][110] = 5'b10000; w[34][111] = 5'b10000; w[34][112] = 5'b10000; w[34][113] = 5'b10000; w[34][114] = 5'b00000; w[34][115] = 5'b10000; w[34][116] = 5'b10000; w[34][117] = 5'b10000; w[34][118] = 5'b00000; w[34][119] = 5'b00000; w[34][120] = 5'b10000; w[34][121] = 5'b10000; w[34][122] = 5'b10000; w[34][123] = 5'b00000; w[34][124] = 5'b10000; w[34][125] = 5'b10000; w[34][126] = 5'b10000; w[34][127] = 5'b10000; w[34][128] = 5'b00000; w[34][129] = 5'b10000; w[34][130] = 5'b10000; w[34][131] = 5'b10000; w[34][132] = 5'b01111; w[34][133] = 5'b00000; w[34][134] = 5'b10000; w[34][135] = 5'b10000; w[34][136] = 5'b10000; w[34][137] = 5'b00000; w[34][138] = 5'b10000; w[34][139] = 5'b10000; w[34][140] = 5'b10000; w[34][141] = 5'b10000; w[34][142] = 5'b00000; w[34][143] = 5'b10000; w[34][144] = 5'b10000; w[34][145] = 5'b10000; w[34][146] = 5'b01111; w[34][147] = 5'b00000; w[34][148] = 5'b10000; w[34][149] = 5'b10000; w[34][150] = 5'b10000; w[34][151] = 5'b00000; w[34][152] = 5'b10000; w[34][153] = 5'b10000; w[34][154] = 5'b10000; w[34][155] = 5'b10000; w[34][156] = 5'b10000; w[34][157] = 5'b10000; w[34][158] = 5'b10000; w[34][159] = 5'b01111; w[34][160] = 5'b01111; w[34][161] = 5'b01111; w[34][162] = 5'b00000; w[34][163] = 5'b10000; w[34][164] = 5'b10000; w[34][165] = 5'b10000; w[34][166] = 5'b10000; w[34][167] = 5'b10000; w[34][168] = 5'b10000; w[34][169] = 5'b10000; w[34][170] = 5'b10000; w[34][171] = 5'b10000; w[34][172] = 5'b10000; w[34][173] = 5'b01111; w[34][174] = 5'b01111; w[34][175] = 5'b01111; w[34][176] = 5'b00000; w[34][177] = 5'b10000; w[34][178] = 5'b10000; w[34][179] = 5'b10000; w[34][180] = 5'b10000; w[34][181] = 5'b10000; w[34][182] = 5'b10000; w[34][183] = 5'b10000; w[34][184] = 5'b10000; w[34][185] = 5'b10000; w[34][186] = 5'b10000; w[34][187] = 5'b10000; w[34][188] = 5'b10000; w[34][189] = 5'b10000; w[34][190] = 5'b10000; w[34][191] = 5'b10000; w[34][192] = 5'b10000; w[34][193] = 5'b10000; w[34][194] = 5'b10000; w[34][195] = 5'b10000; w[34][196] = 5'b10000; w[34][197] = 5'b10000; w[34][198] = 5'b10000; w[34][199] = 5'b10000; w[34][200] = 5'b10000; w[34][201] = 5'b10000; w[34][202] = 5'b10000; w[34][203] = 5'b10000; w[34][204] = 5'b10000; w[34][205] = 5'b10000; w[34][206] = 5'b10000; w[34][207] = 5'b10000; w[34][208] = 5'b10000; w[34][209] = 5'b10000; 
w[35][0] = 5'b10000; w[35][1] = 5'b10000; w[35][2] = 5'b10000; w[35][3] = 5'b10000; w[35][4] = 5'b10000; w[35][5] = 5'b10000; w[35][6] = 5'b10000; w[35][7] = 5'b10000; w[35][8] = 5'b10000; w[35][9] = 5'b10000; w[35][10] = 5'b10000; w[35][11] = 5'b10000; w[35][12] = 5'b10000; w[35][13] = 5'b10000; w[35][14] = 5'b10000; w[35][15] = 5'b10000; w[35][16] = 5'b10000; w[35][17] = 5'b10000; w[35][18] = 5'b10000; w[35][19] = 5'b10000; w[35][20] = 5'b10000; w[35][21] = 5'b10000; w[35][22] = 5'b10000; w[35][23] = 5'b10000; w[35][24] = 5'b10000; w[35][25] = 5'b10000; w[35][26] = 5'b10000; w[35][27] = 5'b10000; w[35][28] = 5'b10000; w[35][29] = 5'b10000; w[35][30] = 5'b00000; w[35][31] = 5'b10000; w[35][32] = 5'b00000; w[35][33] = 5'b01111; w[35][34] = 5'b01111; w[35][35] = 5'b00000; w[35][36] = 5'b01111; w[35][37] = 5'b00000; w[35][38] = 5'b10000; w[35][39] = 5'b00000; w[35][40] = 5'b10000; w[35][41] = 5'b10000; w[35][42] = 5'b10000; w[35][43] = 5'b10000; w[35][44] = 5'b00000; w[35][45] = 5'b00000; w[35][46] = 5'b00000; w[35][47] = 5'b01111; w[35][48] = 5'b01111; w[35][49] = 5'b01111; w[35][50] = 5'b01111; w[35][51] = 5'b00000; w[35][52] = 5'b00000; w[35][53] = 5'b00000; w[35][54] = 5'b10000; w[35][55] = 5'b10000; w[35][56] = 5'b10000; w[35][57] = 5'b10000; w[35][58] = 5'b00000; w[35][59] = 5'b10000; w[35][60] = 5'b10000; w[35][61] = 5'b10000; w[35][62] = 5'b00000; w[35][63] = 5'b01111; w[35][64] = 5'b10000; w[35][65] = 5'b10000; w[35][66] = 5'b10000; w[35][67] = 5'b00000; w[35][68] = 5'b10000; w[35][69] = 5'b10000; w[35][70] = 5'b10000; w[35][71] = 5'b10000; w[35][72] = 5'b00000; w[35][73] = 5'b10000; w[35][74] = 5'b10000; w[35][75] = 5'b10000; w[35][76] = 5'b00000; w[35][77] = 5'b01111; w[35][78] = 5'b10000; w[35][79] = 5'b10000; w[35][80] = 5'b10000; w[35][81] = 5'b00000; w[35][82] = 5'b10000; w[35][83] = 5'b10000; w[35][84] = 5'b10000; w[35][85] = 5'b10000; w[35][86] = 5'b00000; w[35][87] = 5'b10000; w[35][88] = 5'b10000; w[35][89] = 5'b10000; w[35][90] = 5'b00000; w[35][91] = 5'b00000; w[35][92] = 5'b10000; w[35][93] = 5'b10000; w[35][94] = 5'b10000; w[35][95] = 5'b10000; w[35][96] = 5'b10000; w[35][97] = 5'b10000; w[35][98] = 5'b10000; w[35][99] = 5'b10000; w[35][100] = 5'b00000; w[35][101] = 5'b10000; w[35][102] = 5'b10000; w[35][103] = 5'b10000; w[35][104] = 5'b00000; w[35][105] = 5'b00000; w[35][106] = 5'b00000; w[35][107] = 5'b10000; w[35][108] = 5'b10000; w[35][109] = 5'b00000; w[35][110] = 5'b10000; w[35][111] = 5'b10000; w[35][112] = 5'b10000; w[35][113] = 5'b10000; w[35][114] = 5'b00000; w[35][115] = 5'b10000; w[35][116] = 5'b10000; w[35][117] = 5'b10000; w[35][118] = 5'b00000; w[35][119] = 5'b00000; w[35][120] = 5'b10000; w[35][121] = 5'b10000; w[35][122] = 5'b10000; w[35][123] = 5'b00000; w[35][124] = 5'b10000; w[35][125] = 5'b10000; w[35][126] = 5'b10000; w[35][127] = 5'b10000; w[35][128] = 5'b00000; w[35][129] = 5'b10000; w[35][130] = 5'b10000; w[35][131] = 5'b10000; w[35][132] = 5'b01111; w[35][133] = 5'b00000; w[35][134] = 5'b10000; w[35][135] = 5'b10000; w[35][136] = 5'b10000; w[35][137] = 5'b00000; w[35][138] = 5'b10000; w[35][139] = 5'b10000; w[35][140] = 5'b10000; w[35][141] = 5'b10000; w[35][142] = 5'b00000; w[35][143] = 5'b10000; w[35][144] = 5'b10000; w[35][145] = 5'b10000; w[35][146] = 5'b01111; w[35][147] = 5'b00000; w[35][148] = 5'b10000; w[35][149] = 5'b10000; w[35][150] = 5'b10000; w[35][151] = 5'b00000; w[35][152] = 5'b10000; w[35][153] = 5'b10000; w[35][154] = 5'b10000; w[35][155] = 5'b10000; w[35][156] = 5'b10000; w[35][157] = 5'b10000; w[35][158] = 5'b10000; w[35][159] = 5'b01111; w[35][160] = 5'b01111; w[35][161] = 5'b01111; w[35][162] = 5'b00000; w[35][163] = 5'b10000; w[35][164] = 5'b10000; w[35][165] = 5'b10000; w[35][166] = 5'b10000; w[35][167] = 5'b10000; w[35][168] = 5'b10000; w[35][169] = 5'b10000; w[35][170] = 5'b10000; w[35][171] = 5'b10000; w[35][172] = 5'b10000; w[35][173] = 5'b01111; w[35][174] = 5'b01111; w[35][175] = 5'b01111; w[35][176] = 5'b00000; w[35][177] = 5'b10000; w[35][178] = 5'b10000; w[35][179] = 5'b10000; w[35][180] = 5'b10000; w[35][181] = 5'b10000; w[35][182] = 5'b10000; w[35][183] = 5'b10000; w[35][184] = 5'b10000; w[35][185] = 5'b10000; w[35][186] = 5'b10000; w[35][187] = 5'b10000; w[35][188] = 5'b10000; w[35][189] = 5'b10000; w[35][190] = 5'b10000; w[35][191] = 5'b10000; w[35][192] = 5'b10000; w[35][193] = 5'b10000; w[35][194] = 5'b10000; w[35][195] = 5'b10000; w[35][196] = 5'b10000; w[35][197] = 5'b10000; w[35][198] = 5'b10000; w[35][199] = 5'b10000; w[35][200] = 5'b10000; w[35][201] = 5'b10000; w[35][202] = 5'b10000; w[35][203] = 5'b10000; w[35][204] = 5'b10000; w[35][205] = 5'b10000; w[35][206] = 5'b10000; w[35][207] = 5'b10000; w[35][208] = 5'b10000; w[35][209] = 5'b10000; 
w[36][0] = 5'b10000; w[36][1] = 5'b10000; w[36][2] = 5'b10000; w[36][3] = 5'b10000; w[36][4] = 5'b10000; w[36][5] = 5'b10000; w[36][6] = 5'b10000; w[36][7] = 5'b10000; w[36][8] = 5'b10000; w[36][9] = 5'b10000; w[36][10] = 5'b10000; w[36][11] = 5'b10000; w[36][12] = 5'b10000; w[36][13] = 5'b10000; w[36][14] = 5'b10000; w[36][15] = 5'b10000; w[36][16] = 5'b10000; w[36][17] = 5'b10000; w[36][18] = 5'b10000; w[36][19] = 5'b10000; w[36][20] = 5'b10000; w[36][21] = 5'b10000; w[36][22] = 5'b10000; w[36][23] = 5'b10000; w[36][24] = 5'b10000; w[36][25] = 5'b10000; w[36][26] = 5'b10000; w[36][27] = 5'b10000; w[36][28] = 5'b10000; w[36][29] = 5'b10000; w[36][30] = 5'b00000; w[36][31] = 5'b10000; w[36][32] = 5'b00000; w[36][33] = 5'b01111; w[36][34] = 5'b01111; w[36][35] = 5'b01111; w[36][36] = 5'b00000; w[36][37] = 5'b00000; w[36][38] = 5'b10000; w[36][39] = 5'b00000; w[36][40] = 5'b10000; w[36][41] = 5'b10000; w[36][42] = 5'b10000; w[36][43] = 5'b10000; w[36][44] = 5'b00000; w[36][45] = 5'b00000; w[36][46] = 5'b00000; w[36][47] = 5'b01111; w[36][48] = 5'b01111; w[36][49] = 5'b01111; w[36][50] = 5'b01111; w[36][51] = 5'b00000; w[36][52] = 5'b00000; w[36][53] = 5'b00000; w[36][54] = 5'b10000; w[36][55] = 5'b10000; w[36][56] = 5'b10000; w[36][57] = 5'b10000; w[36][58] = 5'b00000; w[36][59] = 5'b10000; w[36][60] = 5'b10000; w[36][61] = 5'b10000; w[36][62] = 5'b00000; w[36][63] = 5'b01111; w[36][64] = 5'b10000; w[36][65] = 5'b10000; w[36][66] = 5'b10000; w[36][67] = 5'b00000; w[36][68] = 5'b10000; w[36][69] = 5'b10000; w[36][70] = 5'b10000; w[36][71] = 5'b10000; w[36][72] = 5'b00000; w[36][73] = 5'b10000; w[36][74] = 5'b10000; w[36][75] = 5'b10000; w[36][76] = 5'b00000; w[36][77] = 5'b01111; w[36][78] = 5'b10000; w[36][79] = 5'b10000; w[36][80] = 5'b10000; w[36][81] = 5'b00000; w[36][82] = 5'b10000; w[36][83] = 5'b10000; w[36][84] = 5'b10000; w[36][85] = 5'b10000; w[36][86] = 5'b00000; w[36][87] = 5'b10000; w[36][88] = 5'b10000; w[36][89] = 5'b10000; w[36][90] = 5'b00000; w[36][91] = 5'b00000; w[36][92] = 5'b10000; w[36][93] = 5'b10000; w[36][94] = 5'b10000; w[36][95] = 5'b10000; w[36][96] = 5'b10000; w[36][97] = 5'b10000; w[36][98] = 5'b10000; w[36][99] = 5'b10000; w[36][100] = 5'b00000; w[36][101] = 5'b10000; w[36][102] = 5'b10000; w[36][103] = 5'b10000; w[36][104] = 5'b00000; w[36][105] = 5'b00000; w[36][106] = 5'b00000; w[36][107] = 5'b10000; w[36][108] = 5'b10000; w[36][109] = 5'b00000; w[36][110] = 5'b10000; w[36][111] = 5'b10000; w[36][112] = 5'b10000; w[36][113] = 5'b10000; w[36][114] = 5'b00000; w[36][115] = 5'b10000; w[36][116] = 5'b10000; w[36][117] = 5'b10000; w[36][118] = 5'b00000; w[36][119] = 5'b00000; w[36][120] = 5'b10000; w[36][121] = 5'b10000; w[36][122] = 5'b10000; w[36][123] = 5'b00000; w[36][124] = 5'b10000; w[36][125] = 5'b10000; w[36][126] = 5'b10000; w[36][127] = 5'b10000; w[36][128] = 5'b00000; w[36][129] = 5'b10000; w[36][130] = 5'b10000; w[36][131] = 5'b10000; w[36][132] = 5'b01111; w[36][133] = 5'b00000; w[36][134] = 5'b10000; w[36][135] = 5'b10000; w[36][136] = 5'b10000; w[36][137] = 5'b00000; w[36][138] = 5'b10000; w[36][139] = 5'b10000; w[36][140] = 5'b10000; w[36][141] = 5'b10000; w[36][142] = 5'b00000; w[36][143] = 5'b10000; w[36][144] = 5'b10000; w[36][145] = 5'b10000; w[36][146] = 5'b01111; w[36][147] = 5'b00000; w[36][148] = 5'b10000; w[36][149] = 5'b10000; w[36][150] = 5'b10000; w[36][151] = 5'b00000; w[36][152] = 5'b10000; w[36][153] = 5'b10000; w[36][154] = 5'b10000; w[36][155] = 5'b10000; w[36][156] = 5'b10000; w[36][157] = 5'b10000; w[36][158] = 5'b10000; w[36][159] = 5'b01111; w[36][160] = 5'b01111; w[36][161] = 5'b01111; w[36][162] = 5'b00000; w[36][163] = 5'b10000; w[36][164] = 5'b10000; w[36][165] = 5'b10000; w[36][166] = 5'b10000; w[36][167] = 5'b10000; w[36][168] = 5'b10000; w[36][169] = 5'b10000; w[36][170] = 5'b10000; w[36][171] = 5'b10000; w[36][172] = 5'b10000; w[36][173] = 5'b01111; w[36][174] = 5'b01111; w[36][175] = 5'b01111; w[36][176] = 5'b00000; w[36][177] = 5'b10000; w[36][178] = 5'b10000; w[36][179] = 5'b10000; w[36][180] = 5'b10000; w[36][181] = 5'b10000; w[36][182] = 5'b10000; w[36][183] = 5'b10000; w[36][184] = 5'b10000; w[36][185] = 5'b10000; w[36][186] = 5'b10000; w[36][187] = 5'b10000; w[36][188] = 5'b10000; w[36][189] = 5'b10000; w[36][190] = 5'b10000; w[36][191] = 5'b10000; w[36][192] = 5'b10000; w[36][193] = 5'b10000; w[36][194] = 5'b10000; w[36][195] = 5'b10000; w[36][196] = 5'b10000; w[36][197] = 5'b10000; w[36][198] = 5'b10000; w[36][199] = 5'b10000; w[36][200] = 5'b10000; w[36][201] = 5'b10000; w[36][202] = 5'b10000; w[36][203] = 5'b10000; w[36][204] = 5'b10000; w[36][205] = 5'b10000; w[36][206] = 5'b10000; w[36][207] = 5'b10000; w[36][208] = 5'b10000; w[36][209] = 5'b10000; 
w[37][0] = 5'b10000; w[37][1] = 5'b10000; w[37][2] = 5'b10000; w[37][3] = 5'b10000; w[37][4] = 5'b10000; w[37][5] = 5'b10000; w[37][6] = 5'b10000; w[37][7] = 5'b10000; w[37][8] = 5'b10000; w[37][9] = 5'b10000; w[37][10] = 5'b10000; w[37][11] = 5'b10000; w[37][12] = 5'b10000; w[37][13] = 5'b10000; w[37][14] = 5'b10000; w[37][15] = 5'b10000; w[37][16] = 5'b10000; w[37][17] = 5'b10000; w[37][18] = 5'b10000; w[37][19] = 5'b10000; w[37][20] = 5'b10000; w[37][21] = 5'b10000; w[37][22] = 5'b10000; w[37][23] = 5'b10000; w[37][24] = 5'b10000; w[37][25] = 5'b10000; w[37][26] = 5'b10000; w[37][27] = 5'b10000; w[37][28] = 5'b10000; w[37][29] = 5'b10000; w[37][30] = 5'b00000; w[37][31] = 5'b01111; w[37][32] = 5'b01111; w[37][33] = 5'b01111; w[37][34] = 5'b00000; w[37][35] = 5'b00000; w[37][36] = 5'b00000; w[37][37] = 5'b00000; w[37][38] = 5'b01111; w[37][39] = 5'b00000; w[37][40] = 5'b10000; w[37][41] = 5'b10000; w[37][42] = 5'b10000; w[37][43] = 5'b10000; w[37][44] = 5'b00000; w[37][45] = 5'b01111; w[37][46] = 5'b01111; w[37][47] = 5'b01111; w[37][48] = 5'b00000; w[37][49] = 5'b00000; w[37][50] = 5'b00000; w[37][51] = 5'b01111; w[37][52] = 5'b01111; w[37][53] = 5'b00000; w[37][54] = 5'b10000; w[37][55] = 5'b10000; w[37][56] = 5'b10000; w[37][57] = 5'b10000; w[37][58] = 5'b00000; w[37][59] = 5'b01111; w[37][60] = 5'b01111; w[37][61] = 5'b00000; w[37][62] = 5'b00000; w[37][63] = 5'b10000; w[37][64] = 5'b10000; w[37][65] = 5'b01111; w[37][66] = 5'b01111; w[37][67] = 5'b00000; w[37][68] = 5'b10000; w[37][69] = 5'b10000; w[37][70] = 5'b10000; w[37][71] = 5'b10000; w[37][72] = 5'b00000; w[37][73] = 5'b01111; w[37][74] = 5'b00000; w[37][75] = 5'b00000; w[37][76] = 5'b00000; w[37][77] = 5'b10000; w[37][78] = 5'b10000; w[37][79] = 5'b00000; w[37][80] = 5'b01111; w[37][81] = 5'b00000; w[37][82] = 5'b10000; w[37][83] = 5'b10000; w[37][84] = 5'b10000; w[37][85] = 5'b10000; w[37][86] = 5'b00000; w[37][87] = 5'b01111; w[37][88] = 5'b00000; w[37][89] = 5'b00000; w[37][90] = 5'b00000; w[37][91] = 5'b00000; w[37][92] = 5'b10000; w[37][93] = 5'b00000; w[37][94] = 5'b00000; w[37][95] = 5'b10000; w[37][96] = 5'b10000; w[37][97] = 5'b10000; w[37][98] = 5'b10000; w[37][99] = 5'b10000; w[37][100] = 5'b00000; w[37][101] = 5'b01111; w[37][102] = 5'b00000; w[37][103] = 5'b10000; w[37][104] = 5'b00000; w[37][105] = 5'b00000; w[37][106] = 5'b00000; w[37][107] = 5'b01111; w[37][108] = 5'b01111; w[37][109] = 5'b00000; w[37][110] = 5'b10000; w[37][111] = 5'b10000; w[37][112] = 5'b10000; w[37][113] = 5'b10000; w[37][114] = 5'b00000; w[37][115] = 5'b01111; w[37][116] = 5'b00000; w[37][117] = 5'b10000; w[37][118] = 5'b00000; w[37][119] = 5'b00000; w[37][120] = 5'b01111; w[37][121] = 5'b01111; w[37][122] = 5'b01111; w[37][123] = 5'b00000; w[37][124] = 5'b10000; w[37][125] = 5'b10000; w[37][126] = 5'b10000; w[37][127] = 5'b10000; w[37][128] = 5'b00000; w[37][129] = 5'b01111; w[37][130] = 5'b00000; w[37][131] = 5'b10000; w[37][132] = 5'b10000; w[37][133] = 5'b00000; w[37][134] = 5'b00000; w[37][135] = 5'b00000; w[37][136] = 5'b01111; w[37][137] = 5'b00000; w[37][138] = 5'b10000; w[37][139] = 5'b10000; w[37][140] = 5'b10000; w[37][141] = 5'b10000; w[37][142] = 5'b00000; w[37][143] = 5'b01111; w[37][144] = 5'b01111; w[37][145] = 5'b10000; w[37][146] = 5'b10000; w[37][147] = 5'b00000; w[37][148] = 5'b00000; w[37][149] = 5'b01111; w[37][150] = 5'b01111; w[37][151] = 5'b00000; w[37][152] = 5'b10000; w[37][153] = 5'b10000; w[37][154] = 5'b10000; w[37][155] = 5'b10000; w[37][156] = 5'b10000; w[37][157] = 5'b01111; w[37][158] = 5'b01111; w[37][159] = 5'b10000; w[37][160] = 5'b00000; w[37][161] = 5'b00000; w[37][162] = 5'b00000; w[37][163] = 5'b01111; w[37][164] = 5'b01111; w[37][165] = 5'b10000; w[37][166] = 5'b10000; w[37][167] = 5'b10000; w[37][168] = 5'b10000; w[37][169] = 5'b10000; w[37][170] = 5'b10000; w[37][171] = 5'b00000; w[37][172] = 5'b01111; w[37][173] = 5'b10000; w[37][174] = 5'b00000; w[37][175] = 5'b00000; w[37][176] = 5'b00000; w[37][177] = 5'b01111; w[37][178] = 5'b00000; w[37][179] = 5'b10000; w[37][180] = 5'b10000; w[37][181] = 5'b10000; w[37][182] = 5'b10000; w[37][183] = 5'b10000; w[37][184] = 5'b10000; w[37][185] = 5'b10000; w[37][186] = 5'b10000; w[37][187] = 5'b10000; w[37][188] = 5'b10000; w[37][189] = 5'b10000; w[37][190] = 5'b10000; w[37][191] = 5'b10000; w[37][192] = 5'b10000; w[37][193] = 5'b10000; w[37][194] = 5'b10000; w[37][195] = 5'b10000; w[37][196] = 5'b10000; w[37][197] = 5'b10000; w[37][198] = 5'b10000; w[37][199] = 5'b10000; w[37][200] = 5'b10000; w[37][201] = 5'b10000; w[37][202] = 5'b10000; w[37][203] = 5'b10000; w[37][204] = 5'b10000; w[37][205] = 5'b10000; w[37][206] = 5'b10000; w[37][207] = 5'b10000; w[37][208] = 5'b10000; w[37][209] = 5'b10000; 
w[38][0] = 5'b00000; w[38][1] = 5'b00000; w[38][2] = 5'b00000; w[38][3] = 5'b00000; w[38][4] = 5'b00000; w[38][5] = 5'b00000; w[38][6] = 5'b00000; w[38][7] = 5'b00000; w[38][8] = 5'b00000; w[38][9] = 5'b00000; w[38][10] = 5'b00000; w[38][11] = 5'b00000; w[38][12] = 5'b00000; w[38][13] = 5'b00000; w[38][14] = 5'b00000; w[38][15] = 5'b00000; w[38][16] = 5'b00000; w[38][17] = 5'b00000; w[38][18] = 5'b00000; w[38][19] = 5'b00000; w[38][20] = 5'b00000; w[38][21] = 5'b00000; w[38][22] = 5'b00000; w[38][23] = 5'b00000; w[38][24] = 5'b00000; w[38][25] = 5'b00000; w[38][26] = 5'b00000; w[38][27] = 5'b00000; w[38][28] = 5'b00000; w[38][29] = 5'b00000; w[38][30] = 5'b01111; w[38][31] = 5'b01111; w[38][32] = 5'b01111; w[38][33] = 5'b00000; w[38][34] = 5'b10000; w[38][35] = 5'b10000; w[38][36] = 5'b10000; w[38][37] = 5'b01111; w[38][38] = 5'b00000; w[38][39] = 5'b01111; w[38][40] = 5'b00000; w[38][41] = 5'b00000; w[38][42] = 5'b00000; w[38][43] = 5'b00000; w[38][44] = 5'b01111; w[38][45] = 5'b01111; w[38][46] = 5'b01111; w[38][47] = 5'b00000; w[38][48] = 5'b10000; w[38][49] = 5'b10000; w[38][50] = 5'b10000; w[38][51] = 5'b01111; w[38][52] = 5'b01111; w[38][53] = 5'b01111; w[38][54] = 5'b00000; w[38][55] = 5'b00000; w[38][56] = 5'b00000; w[38][57] = 5'b00000; w[38][58] = 5'b10000; w[38][59] = 5'b00000; w[38][60] = 5'b00000; w[38][61] = 5'b01111; w[38][62] = 5'b01111; w[38][63] = 5'b00000; w[38][64] = 5'b00000; w[38][65] = 5'b00000; w[38][66] = 5'b00000; w[38][67] = 5'b10000; w[38][68] = 5'b00000; w[38][69] = 5'b00000; w[38][70] = 5'b00000; w[38][71] = 5'b00000; w[38][72] = 5'b10000; w[38][73] = 5'b00000; w[38][74] = 5'b01111; w[38][75] = 5'b01111; w[38][76] = 5'b01111; w[38][77] = 5'b00000; w[38][78] = 5'b00000; w[38][79] = 5'b01111; w[38][80] = 5'b00000; w[38][81] = 5'b10000; w[38][82] = 5'b00000; w[38][83] = 5'b00000; w[38][84] = 5'b00000; w[38][85] = 5'b00000; w[38][86] = 5'b10000; w[38][87] = 5'b00000; w[38][88] = 5'b01111; w[38][89] = 5'b01111; w[38][90] = 5'b01111; w[38][91] = 5'b01111; w[38][92] = 5'b00000; w[38][93] = 5'b01111; w[38][94] = 5'b01111; w[38][95] = 5'b00000; w[38][96] = 5'b00000; w[38][97] = 5'b00000; w[38][98] = 5'b00000; w[38][99] = 5'b00000; w[38][100] = 5'b10000; w[38][101] = 5'b00000; w[38][102] = 5'b01111; w[38][103] = 5'b00000; w[38][104] = 5'b01111; w[38][105] = 5'b01111; w[38][106] = 5'b10000; w[38][107] = 5'b00000; w[38][108] = 5'b00000; w[38][109] = 5'b10000; w[38][110] = 5'b00000; w[38][111] = 5'b00000; w[38][112] = 5'b00000; w[38][113] = 5'b00000; w[38][114] = 5'b10000; w[38][115] = 5'b00000; w[38][116] = 5'b01111; w[38][117] = 5'b00000; w[38][118] = 5'b01111; w[38][119] = 5'b01111; w[38][120] = 5'b00000; w[38][121] = 5'b00000; w[38][122] = 5'b00000; w[38][123] = 5'b10000; w[38][124] = 5'b00000; w[38][125] = 5'b00000; w[38][126] = 5'b00000; w[38][127] = 5'b00000; w[38][128] = 5'b10000; w[38][129] = 5'b00000; w[38][130] = 5'b01111; w[38][131] = 5'b00000; w[38][132] = 5'b00000; w[38][133] = 5'b01111; w[38][134] = 5'b01111; w[38][135] = 5'b01111; w[38][136] = 5'b00000; w[38][137] = 5'b10000; w[38][138] = 5'b00000; w[38][139] = 5'b00000; w[38][140] = 5'b00000; w[38][141] = 5'b00000; w[38][142] = 5'b10000; w[38][143] = 5'b00000; w[38][144] = 5'b00000; w[38][145] = 5'b00000; w[38][146] = 5'b00000; w[38][147] = 5'b01111; w[38][148] = 5'b01111; w[38][149] = 5'b00000; w[38][150] = 5'b00000; w[38][151] = 5'b10000; w[38][152] = 5'b00000; w[38][153] = 5'b00000; w[38][154] = 5'b00000; w[38][155] = 5'b00000; w[38][156] = 5'b00000; w[38][157] = 5'b00000; w[38][158] = 5'b00000; w[38][159] = 5'b10000; w[38][160] = 5'b10000; w[38][161] = 5'b10000; w[38][162] = 5'b10000; w[38][163] = 5'b00000; w[38][164] = 5'b00000; w[38][165] = 5'b00000; w[38][166] = 5'b00000; w[38][167] = 5'b00000; w[38][168] = 5'b00000; w[38][169] = 5'b00000; w[38][170] = 5'b00000; w[38][171] = 5'b01111; w[38][172] = 5'b00000; w[38][173] = 5'b10000; w[38][174] = 5'b10000; w[38][175] = 5'b10000; w[38][176] = 5'b10000; w[38][177] = 5'b00000; w[38][178] = 5'b01111; w[38][179] = 5'b00000; w[38][180] = 5'b00000; w[38][181] = 5'b00000; w[38][182] = 5'b00000; w[38][183] = 5'b00000; w[38][184] = 5'b00000; w[38][185] = 5'b00000; w[38][186] = 5'b00000; w[38][187] = 5'b00000; w[38][188] = 5'b00000; w[38][189] = 5'b00000; w[38][190] = 5'b00000; w[38][191] = 5'b00000; w[38][192] = 5'b00000; w[38][193] = 5'b00000; w[38][194] = 5'b00000; w[38][195] = 5'b00000; w[38][196] = 5'b00000; w[38][197] = 5'b00000; w[38][198] = 5'b00000; w[38][199] = 5'b00000; w[38][200] = 5'b00000; w[38][201] = 5'b00000; w[38][202] = 5'b00000; w[38][203] = 5'b00000; w[38][204] = 5'b00000; w[38][205] = 5'b00000; w[38][206] = 5'b00000; w[38][207] = 5'b00000; w[38][208] = 5'b00000; w[38][209] = 5'b00000; 
w[39][0] = 5'b01111; w[39][1] = 5'b01111; w[39][2] = 5'b01111; w[39][3] = 5'b01111; w[39][4] = 5'b01111; w[39][5] = 5'b01111; w[39][6] = 5'b01111; w[39][7] = 5'b01111; w[39][8] = 5'b01111; w[39][9] = 5'b01111; w[39][10] = 5'b01111; w[39][11] = 5'b01111; w[39][12] = 5'b01111; w[39][13] = 5'b01111; w[39][14] = 5'b01111; w[39][15] = 5'b01111; w[39][16] = 5'b01111; w[39][17] = 5'b01111; w[39][18] = 5'b01111; w[39][19] = 5'b01111; w[39][20] = 5'b01111; w[39][21] = 5'b01111; w[39][22] = 5'b01111; w[39][23] = 5'b01111; w[39][24] = 5'b01111; w[39][25] = 5'b01111; w[39][26] = 5'b01111; w[39][27] = 5'b01111; w[39][28] = 5'b01111; w[39][29] = 5'b01111; w[39][30] = 5'b01111; w[39][31] = 5'b01111; w[39][32] = 5'b00000; w[39][33] = 5'b10000; w[39][34] = 5'b00000; w[39][35] = 5'b00000; w[39][36] = 5'b00000; w[39][37] = 5'b00000; w[39][38] = 5'b01111; w[39][39] = 5'b00000; w[39][40] = 5'b01111; w[39][41] = 5'b01111; w[39][42] = 5'b01111; w[39][43] = 5'b01111; w[39][44] = 5'b01111; w[39][45] = 5'b00000; w[39][46] = 5'b00000; w[39][47] = 5'b10000; w[39][48] = 5'b00000; w[39][49] = 5'b00000; w[39][50] = 5'b00000; w[39][51] = 5'b00000; w[39][52] = 5'b00000; w[39][53] = 5'b01111; w[39][54] = 5'b01111; w[39][55] = 5'b01111; w[39][56] = 5'b01111; w[39][57] = 5'b01111; w[39][58] = 5'b00000; w[39][59] = 5'b10000; w[39][60] = 5'b10000; w[39][61] = 5'b00000; w[39][62] = 5'b00000; w[39][63] = 5'b01111; w[39][64] = 5'b01111; w[39][65] = 5'b10000; w[39][66] = 5'b10000; w[39][67] = 5'b00000; w[39][68] = 5'b01111; w[39][69] = 5'b01111; w[39][70] = 5'b01111; w[39][71] = 5'b01111; w[39][72] = 5'b00000; w[39][73] = 5'b10000; w[39][74] = 5'b00000; w[39][75] = 5'b00000; w[39][76] = 5'b00000; w[39][77] = 5'b01111; w[39][78] = 5'b01111; w[39][79] = 5'b00000; w[39][80] = 5'b10000; w[39][81] = 5'b00000; w[39][82] = 5'b01111; w[39][83] = 5'b01111; w[39][84] = 5'b01111; w[39][85] = 5'b01111; w[39][86] = 5'b00000; w[39][87] = 5'b10000; w[39][88] = 5'b00000; w[39][89] = 5'b00000; w[39][90] = 5'b00000; w[39][91] = 5'b00000; w[39][92] = 5'b01111; w[39][93] = 5'b00000; w[39][94] = 5'b00000; w[39][95] = 5'b01111; w[39][96] = 5'b01111; w[39][97] = 5'b01111; w[39][98] = 5'b01111; w[39][99] = 5'b01111; w[39][100] = 5'b00000; w[39][101] = 5'b10000; w[39][102] = 5'b00000; w[39][103] = 5'b01111; w[39][104] = 5'b00000; w[39][105] = 5'b00000; w[39][106] = 5'b00000; w[39][107] = 5'b10000; w[39][108] = 5'b10000; w[39][109] = 5'b00000; w[39][110] = 5'b01111; w[39][111] = 5'b01111; w[39][112] = 5'b01111; w[39][113] = 5'b01111; w[39][114] = 5'b00000; w[39][115] = 5'b10000; w[39][116] = 5'b00000; w[39][117] = 5'b01111; w[39][118] = 5'b00000; w[39][119] = 5'b00000; w[39][120] = 5'b10000; w[39][121] = 5'b10000; w[39][122] = 5'b10000; w[39][123] = 5'b00000; w[39][124] = 5'b01111; w[39][125] = 5'b01111; w[39][126] = 5'b01111; w[39][127] = 5'b01111; w[39][128] = 5'b00000; w[39][129] = 5'b10000; w[39][130] = 5'b00000; w[39][131] = 5'b01111; w[39][132] = 5'b01111; w[39][133] = 5'b00000; w[39][134] = 5'b00000; w[39][135] = 5'b00000; w[39][136] = 5'b10000; w[39][137] = 5'b00000; w[39][138] = 5'b01111; w[39][139] = 5'b01111; w[39][140] = 5'b01111; w[39][141] = 5'b01111; w[39][142] = 5'b00000; w[39][143] = 5'b10000; w[39][144] = 5'b10000; w[39][145] = 5'b01111; w[39][146] = 5'b01111; w[39][147] = 5'b00000; w[39][148] = 5'b00000; w[39][149] = 5'b10000; w[39][150] = 5'b10000; w[39][151] = 5'b00000; w[39][152] = 5'b01111; w[39][153] = 5'b01111; w[39][154] = 5'b01111; w[39][155] = 5'b01111; w[39][156] = 5'b01111; w[39][157] = 5'b10000; w[39][158] = 5'b10000; w[39][159] = 5'b10000; w[39][160] = 5'b00000; w[39][161] = 5'b00000; w[39][162] = 5'b10000; w[39][163] = 5'b10000; w[39][164] = 5'b10000; w[39][165] = 5'b01111; w[39][166] = 5'b01111; w[39][167] = 5'b01111; w[39][168] = 5'b01111; w[39][169] = 5'b01111; w[39][170] = 5'b01111; w[39][171] = 5'b00000; w[39][172] = 5'b10000; w[39][173] = 5'b10000; w[39][174] = 5'b00000; w[39][175] = 5'b00000; w[39][176] = 5'b10000; w[39][177] = 5'b10000; w[39][178] = 5'b00000; w[39][179] = 5'b01111; w[39][180] = 5'b01111; w[39][181] = 5'b01111; w[39][182] = 5'b01111; w[39][183] = 5'b01111; w[39][184] = 5'b01111; w[39][185] = 5'b01111; w[39][186] = 5'b01111; w[39][187] = 5'b01111; w[39][188] = 5'b01111; w[39][189] = 5'b01111; w[39][190] = 5'b01111; w[39][191] = 5'b01111; w[39][192] = 5'b01111; w[39][193] = 5'b01111; w[39][194] = 5'b01111; w[39][195] = 5'b01111; w[39][196] = 5'b01111; w[39][197] = 5'b01111; w[39][198] = 5'b01111; w[39][199] = 5'b01111; w[39][200] = 5'b01111; w[39][201] = 5'b01111; w[39][202] = 5'b01111; w[39][203] = 5'b01111; w[39][204] = 5'b01111; w[39][205] = 5'b01111; w[39][206] = 5'b01111; w[39][207] = 5'b01111; w[39][208] = 5'b01111; w[39][209] = 5'b01111; 
w[40][0] = 5'b01111; w[40][1] = 5'b01111; w[40][2] = 5'b01111; w[40][3] = 5'b01111; w[40][4] = 5'b01111; w[40][5] = 5'b01111; w[40][6] = 5'b01111; w[40][7] = 5'b01111; w[40][8] = 5'b01111; w[40][9] = 5'b01111; w[40][10] = 5'b01111; w[40][11] = 5'b01111; w[40][12] = 5'b01111; w[40][13] = 5'b01111; w[40][14] = 5'b01111; w[40][15] = 5'b01111; w[40][16] = 5'b01111; w[40][17] = 5'b01111; w[40][18] = 5'b01111; w[40][19] = 5'b01111; w[40][20] = 5'b01111; w[40][21] = 5'b01111; w[40][22] = 5'b01111; w[40][23] = 5'b01111; w[40][24] = 5'b01111; w[40][25] = 5'b01111; w[40][26] = 5'b01111; w[40][27] = 5'b01111; w[40][28] = 5'b01111; w[40][29] = 5'b01111; w[40][30] = 5'b01111; w[40][31] = 5'b00000; w[40][32] = 5'b10000; w[40][33] = 5'b10000; w[40][34] = 5'b10000; w[40][35] = 5'b10000; w[40][36] = 5'b10000; w[40][37] = 5'b10000; w[40][38] = 5'b00000; w[40][39] = 5'b01111; w[40][40] = 5'b00000; w[40][41] = 5'b01111; w[40][42] = 5'b01111; w[40][43] = 5'b01111; w[40][44] = 5'b01111; w[40][45] = 5'b10000; w[40][46] = 5'b10000; w[40][47] = 5'b10000; w[40][48] = 5'b10000; w[40][49] = 5'b10000; w[40][50] = 5'b10000; w[40][51] = 5'b10000; w[40][52] = 5'b10000; w[40][53] = 5'b01111; w[40][54] = 5'b01111; w[40][55] = 5'b01111; w[40][56] = 5'b01111; w[40][57] = 5'b01111; w[40][58] = 5'b01111; w[40][59] = 5'b00000; w[40][60] = 5'b00000; w[40][61] = 5'b01111; w[40][62] = 5'b10000; w[40][63] = 5'b00000; w[40][64] = 5'b01111; w[40][65] = 5'b00000; w[40][66] = 5'b00000; w[40][67] = 5'b01111; w[40][68] = 5'b01111; w[40][69] = 5'b01111; w[40][70] = 5'b01111; w[40][71] = 5'b01111; w[40][72] = 5'b01111; w[40][73] = 5'b00000; w[40][74] = 5'b01111; w[40][75] = 5'b01111; w[40][76] = 5'b10000; w[40][77] = 5'b00000; w[40][78] = 5'b01111; w[40][79] = 5'b01111; w[40][80] = 5'b00000; w[40][81] = 5'b01111; w[40][82] = 5'b01111; w[40][83] = 5'b01111; w[40][84] = 5'b01111; w[40][85] = 5'b01111; w[40][86] = 5'b01111; w[40][87] = 5'b00000; w[40][88] = 5'b01111; w[40][89] = 5'b01111; w[40][90] = 5'b10000; w[40][91] = 5'b10000; w[40][92] = 5'b01111; w[40][93] = 5'b01111; w[40][94] = 5'b01111; w[40][95] = 5'b01111; w[40][96] = 5'b01111; w[40][97] = 5'b01111; w[40][98] = 5'b01111; w[40][99] = 5'b01111; w[40][100] = 5'b01111; w[40][101] = 5'b00000; w[40][102] = 5'b01111; w[40][103] = 5'b01111; w[40][104] = 5'b10000; w[40][105] = 5'b10000; w[40][106] = 5'b01111; w[40][107] = 5'b00000; w[40][108] = 5'b00000; w[40][109] = 5'b01111; w[40][110] = 5'b01111; w[40][111] = 5'b01111; w[40][112] = 5'b01111; w[40][113] = 5'b01111; w[40][114] = 5'b01111; w[40][115] = 5'b00000; w[40][116] = 5'b01111; w[40][117] = 5'b01111; w[40][118] = 5'b10000; w[40][119] = 5'b10000; w[40][120] = 5'b00000; w[40][121] = 5'b00000; w[40][122] = 5'b00000; w[40][123] = 5'b01111; w[40][124] = 5'b01111; w[40][125] = 5'b01111; w[40][126] = 5'b01111; w[40][127] = 5'b01111; w[40][128] = 5'b01111; w[40][129] = 5'b00000; w[40][130] = 5'b01111; w[40][131] = 5'b01111; w[40][132] = 5'b00000; w[40][133] = 5'b10000; w[40][134] = 5'b01111; w[40][135] = 5'b01111; w[40][136] = 5'b00000; w[40][137] = 5'b01111; w[40][138] = 5'b01111; w[40][139] = 5'b01111; w[40][140] = 5'b01111; w[40][141] = 5'b01111; w[40][142] = 5'b01111; w[40][143] = 5'b00000; w[40][144] = 5'b00000; w[40][145] = 5'b01111; w[40][146] = 5'b00000; w[40][147] = 5'b10000; w[40][148] = 5'b01111; w[40][149] = 5'b00000; w[40][150] = 5'b00000; w[40][151] = 5'b01111; w[40][152] = 5'b01111; w[40][153] = 5'b01111; w[40][154] = 5'b01111; w[40][155] = 5'b01111; w[40][156] = 5'b01111; w[40][157] = 5'b00000; w[40][158] = 5'b00000; w[40][159] = 5'b00000; w[40][160] = 5'b10000; w[40][161] = 5'b10000; w[40][162] = 5'b10000; w[40][163] = 5'b00000; w[40][164] = 5'b00000; w[40][165] = 5'b01111; w[40][166] = 5'b01111; w[40][167] = 5'b01111; w[40][168] = 5'b01111; w[40][169] = 5'b01111; w[40][170] = 5'b01111; w[40][171] = 5'b01111; w[40][172] = 5'b00000; w[40][173] = 5'b00000; w[40][174] = 5'b10000; w[40][175] = 5'b10000; w[40][176] = 5'b10000; w[40][177] = 5'b00000; w[40][178] = 5'b01111; w[40][179] = 5'b01111; w[40][180] = 5'b01111; w[40][181] = 5'b01111; w[40][182] = 5'b01111; w[40][183] = 5'b01111; w[40][184] = 5'b01111; w[40][185] = 5'b01111; w[40][186] = 5'b01111; w[40][187] = 5'b01111; w[40][188] = 5'b01111; w[40][189] = 5'b01111; w[40][190] = 5'b01111; w[40][191] = 5'b01111; w[40][192] = 5'b01111; w[40][193] = 5'b01111; w[40][194] = 5'b01111; w[40][195] = 5'b01111; w[40][196] = 5'b01111; w[40][197] = 5'b01111; w[40][198] = 5'b01111; w[40][199] = 5'b01111; w[40][200] = 5'b01111; w[40][201] = 5'b01111; w[40][202] = 5'b01111; w[40][203] = 5'b01111; w[40][204] = 5'b01111; w[40][205] = 5'b01111; w[40][206] = 5'b01111; w[40][207] = 5'b01111; w[40][208] = 5'b01111; w[40][209] = 5'b01111; 
w[41][0] = 5'b01111; w[41][1] = 5'b01111; w[41][2] = 5'b01111; w[41][3] = 5'b01111; w[41][4] = 5'b01111; w[41][5] = 5'b01111; w[41][6] = 5'b01111; w[41][7] = 5'b01111; w[41][8] = 5'b01111; w[41][9] = 5'b01111; w[41][10] = 5'b01111; w[41][11] = 5'b01111; w[41][12] = 5'b01111; w[41][13] = 5'b01111; w[41][14] = 5'b01111; w[41][15] = 5'b01111; w[41][16] = 5'b01111; w[41][17] = 5'b01111; w[41][18] = 5'b01111; w[41][19] = 5'b01111; w[41][20] = 5'b01111; w[41][21] = 5'b01111; w[41][22] = 5'b01111; w[41][23] = 5'b01111; w[41][24] = 5'b01111; w[41][25] = 5'b01111; w[41][26] = 5'b01111; w[41][27] = 5'b01111; w[41][28] = 5'b01111; w[41][29] = 5'b01111; w[41][30] = 5'b01111; w[41][31] = 5'b00000; w[41][32] = 5'b10000; w[41][33] = 5'b10000; w[41][34] = 5'b10000; w[41][35] = 5'b10000; w[41][36] = 5'b10000; w[41][37] = 5'b10000; w[41][38] = 5'b00000; w[41][39] = 5'b01111; w[41][40] = 5'b01111; w[41][41] = 5'b00000; w[41][42] = 5'b01111; w[41][43] = 5'b01111; w[41][44] = 5'b01111; w[41][45] = 5'b10000; w[41][46] = 5'b10000; w[41][47] = 5'b10000; w[41][48] = 5'b10000; w[41][49] = 5'b10000; w[41][50] = 5'b10000; w[41][51] = 5'b10000; w[41][52] = 5'b10000; w[41][53] = 5'b01111; w[41][54] = 5'b01111; w[41][55] = 5'b01111; w[41][56] = 5'b01111; w[41][57] = 5'b01111; w[41][58] = 5'b01111; w[41][59] = 5'b00000; w[41][60] = 5'b00000; w[41][61] = 5'b01111; w[41][62] = 5'b10000; w[41][63] = 5'b00000; w[41][64] = 5'b01111; w[41][65] = 5'b00000; w[41][66] = 5'b00000; w[41][67] = 5'b01111; w[41][68] = 5'b01111; w[41][69] = 5'b01111; w[41][70] = 5'b01111; w[41][71] = 5'b01111; w[41][72] = 5'b01111; w[41][73] = 5'b00000; w[41][74] = 5'b01111; w[41][75] = 5'b01111; w[41][76] = 5'b10000; w[41][77] = 5'b00000; w[41][78] = 5'b01111; w[41][79] = 5'b01111; w[41][80] = 5'b00000; w[41][81] = 5'b01111; w[41][82] = 5'b01111; w[41][83] = 5'b01111; w[41][84] = 5'b01111; w[41][85] = 5'b01111; w[41][86] = 5'b01111; w[41][87] = 5'b00000; w[41][88] = 5'b01111; w[41][89] = 5'b01111; w[41][90] = 5'b10000; w[41][91] = 5'b10000; w[41][92] = 5'b01111; w[41][93] = 5'b01111; w[41][94] = 5'b01111; w[41][95] = 5'b01111; w[41][96] = 5'b01111; w[41][97] = 5'b01111; w[41][98] = 5'b01111; w[41][99] = 5'b01111; w[41][100] = 5'b01111; w[41][101] = 5'b00000; w[41][102] = 5'b01111; w[41][103] = 5'b01111; w[41][104] = 5'b10000; w[41][105] = 5'b10000; w[41][106] = 5'b01111; w[41][107] = 5'b00000; w[41][108] = 5'b00000; w[41][109] = 5'b01111; w[41][110] = 5'b01111; w[41][111] = 5'b01111; w[41][112] = 5'b01111; w[41][113] = 5'b01111; w[41][114] = 5'b01111; w[41][115] = 5'b00000; w[41][116] = 5'b01111; w[41][117] = 5'b01111; w[41][118] = 5'b10000; w[41][119] = 5'b10000; w[41][120] = 5'b00000; w[41][121] = 5'b00000; w[41][122] = 5'b00000; w[41][123] = 5'b01111; w[41][124] = 5'b01111; w[41][125] = 5'b01111; w[41][126] = 5'b01111; w[41][127] = 5'b01111; w[41][128] = 5'b01111; w[41][129] = 5'b00000; w[41][130] = 5'b01111; w[41][131] = 5'b01111; w[41][132] = 5'b00000; w[41][133] = 5'b10000; w[41][134] = 5'b01111; w[41][135] = 5'b01111; w[41][136] = 5'b00000; w[41][137] = 5'b01111; w[41][138] = 5'b01111; w[41][139] = 5'b01111; w[41][140] = 5'b01111; w[41][141] = 5'b01111; w[41][142] = 5'b01111; w[41][143] = 5'b00000; w[41][144] = 5'b00000; w[41][145] = 5'b01111; w[41][146] = 5'b00000; w[41][147] = 5'b10000; w[41][148] = 5'b01111; w[41][149] = 5'b00000; w[41][150] = 5'b00000; w[41][151] = 5'b01111; w[41][152] = 5'b01111; w[41][153] = 5'b01111; w[41][154] = 5'b01111; w[41][155] = 5'b01111; w[41][156] = 5'b01111; w[41][157] = 5'b00000; w[41][158] = 5'b00000; w[41][159] = 5'b00000; w[41][160] = 5'b10000; w[41][161] = 5'b10000; w[41][162] = 5'b10000; w[41][163] = 5'b00000; w[41][164] = 5'b00000; w[41][165] = 5'b01111; w[41][166] = 5'b01111; w[41][167] = 5'b01111; w[41][168] = 5'b01111; w[41][169] = 5'b01111; w[41][170] = 5'b01111; w[41][171] = 5'b01111; w[41][172] = 5'b00000; w[41][173] = 5'b00000; w[41][174] = 5'b10000; w[41][175] = 5'b10000; w[41][176] = 5'b10000; w[41][177] = 5'b00000; w[41][178] = 5'b01111; w[41][179] = 5'b01111; w[41][180] = 5'b01111; w[41][181] = 5'b01111; w[41][182] = 5'b01111; w[41][183] = 5'b01111; w[41][184] = 5'b01111; w[41][185] = 5'b01111; w[41][186] = 5'b01111; w[41][187] = 5'b01111; w[41][188] = 5'b01111; w[41][189] = 5'b01111; w[41][190] = 5'b01111; w[41][191] = 5'b01111; w[41][192] = 5'b01111; w[41][193] = 5'b01111; w[41][194] = 5'b01111; w[41][195] = 5'b01111; w[41][196] = 5'b01111; w[41][197] = 5'b01111; w[41][198] = 5'b01111; w[41][199] = 5'b01111; w[41][200] = 5'b01111; w[41][201] = 5'b01111; w[41][202] = 5'b01111; w[41][203] = 5'b01111; w[41][204] = 5'b01111; w[41][205] = 5'b01111; w[41][206] = 5'b01111; w[41][207] = 5'b01111; w[41][208] = 5'b01111; w[41][209] = 5'b01111; 
w[42][0] = 5'b01111; w[42][1] = 5'b01111; w[42][2] = 5'b01111; w[42][3] = 5'b01111; w[42][4] = 5'b01111; w[42][5] = 5'b01111; w[42][6] = 5'b01111; w[42][7] = 5'b01111; w[42][8] = 5'b01111; w[42][9] = 5'b01111; w[42][10] = 5'b01111; w[42][11] = 5'b01111; w[42][12] = 5'b01111; w[42][13] = 5'b01111; w[42][14] = 5'b01111; w[42][15] = 5'b01111; w[42][16] = 5'b01111; w[42][17] = 5'b01111; w[42][18] = 5'b01111; w[42][19] = 5'b01111; w[42][20] = 5'b01111; w[42][21] = 5'b01111; w[42][22] = 5'b01111; w[42][23] = 5'b01111; w[42][24] = 5'b01111; w[42][25] = 5'b01111; w[42][26] = 5'b01111; w[42][27] = 5'b01111; w[42][28] = 5'b01111; w[42][29] = 5'b01111; w[42][30] = 5'b01111; w[42][31] = 5'b00000; w[42][32] = 5'b10000; w[42][33] = 5'b10000; w[42][34] = 5'b10000; w[42][35] = 5'b10000; w[42][36] = 5'b10000; w[42][37] = 5'b10000; w[42][38] = 5'b00000; w[42][39] = 5'b01111; w[42][40] = 5'b01111; w[42][41] = 5'b01111; w[42][42] = 5'b00000; w[42][43] = 5'b01111; w[42][44] = 5'b01111; w[42][45] = 5'b10000; w[42][46] = 5'b10000; w[42][47] = 5'b10000; w[42][48] = 5'b10000; w[42][49] = 5'b10000; w[42][50] = 5'b10000; w[42][51] = 5'b10000; w[42][52] = 5'b10000; w[42][53] = 5'b01111; w[42][54] = 5'b01111; w[42][55] = 5'b01111; w[42][56] = 5'b01111; w[42][57] = 5'b01111; w[42][58] = 5'b01111; w[42][59] = 5'b00000; w[42][60] = 5'b00000; w[42][61] = 5'b01111; w[42][62] = 5'b10000; w[42][63] = 5'b00000; w[42][64] = 5'b01111; w[42][65] = 5'b00000; w[42][66] = 5'b00000; w[42][67] = 5'b01111; w[42][68] = 5'b01111; w[42][69] = 5'b01111; w[42][70] = 5'b01111; w[42][71] = 5'b01111; w[42][72] = 5'b01111; w[42][73] = 5'b00000; w[42][74] = 5'b01111; w[42][75] = 5'b01111; w[42][76] = 5'b10000; w[42][77] = 5'b00000; w[42][78] = 5'b01111; w[42][79] = 5'b01111; w[42][80] = 5'b00000; w[42][81] = 5'b01111; w[42][82] = 5'b01111; w[42][83] = 5'b01111; w[42][84] = 5'b01111; w[42][85] = 5'b01111; w[42][86] = 5'b01111; w[42][87] = 5'b00000; w[42][88] = 5'b01111; w[42][89] = 5'b01111; w[42][90] = 5'b10000; w[42][91] = 5'b10000; w[42][92] = 5'b01111; w[42][93] = 5'b01111; w[42][94] = 5'b01111; w[42][95] = 5'b01111; w[42][96] = 5'b01111; w[42][97] = 5'b01111; w[42][98] = 5'b01111; w[42][99] = 5'b01111; w[42][100] = 5'b01111; w[42][101] = 5'b00000; w[42][102] = 5'b01111; w[42][103] = 5'b01111; w[42][104] = 5'b10000; w[42][105] = 5'b10000; w[42][106] = 5'b01111; w[42][107] = 5'b00000; w[42][108] = 5'b00000; w[42][109] = 5'b01111; w[42][110] = 5'b01111; w[42][111] = 5'b01111; w[42][112] = 5'b01111; w[42][113] = 5'b01111; w[42][114] = 5'b01111; w[42][115] = 5'b00000; w[42][116] = 5'b01111; w[42][117] = 5'b01111; w[42][118] = 5'b10000; w[42][119] = 5'b10000; w[42][120] = 5'b00000; w[42][121] = 5'b00000; w[42][122] = 5'b00000; w[42][123] = 5'b01111; w[42][124] = 5'b01111; w[42][125] = 5'b01111; w[42][126] = 5'b01111; w[42][127] = 5'b01111; w[42][128] = 5'b01111; w[42][129] = 5'b00000; w[42][130] = 5'b01111; w[42][131] = 5'b01111; w[42][132] = 5'b00000; w[42][133] = 5'b10000; w[42][134] = 5'b01111; w[42][135] = 5'b01111; w[42][136] = 5'b00000; w[42][137] = 5'b01111; w[42][138] = 5'b01111; w[42][139] = 5'b01111; w[42][140] = 5'b01111; w[42][141] = 5'b01111; w[42][142] = 5'b01111; w[42][143] = 5'b00000; w[42][144] = 5'b00000; w[42][145] = 5'b01111; w[42][146] = 5'b00000; w[42][147] = 5'b10000; w[42][148] = 5'b01111; w[42][149] = 5'b00000; w[42][150] = 5'b00000; w[42][151] = 5'b01111; w[42][152] = 5'b01111; w[42][153] = 5'b01111; w[42][154] = 5'b01111; w[42][155] = 5'b01111; w[42][156] = 5'b01111; w[42][157] = 5'b00000; w[42][158] = 5'b00000; w[42][159] = 5'b00000; w[42][160] = 5'b10000; w[42][161] = 5'b10000; w[42][162] = 5'b10000; w[42][163] = 5'b00000; w[42][164] = 5'b00000; w[42][165] = 5'b01111; w[42][166] = 5'b01111; w[42][167] = 5'b01111; w[42][168] = 5'b01111; w[42][169] = 5'b01111; w[42][170] = 5'b01111; w[42][171] = 5'b01111; w[42][172] = 5'b00000; w[42][173] = 5'b00000; w[42][174] = 5'b10000; w[42][175] = 5'b10000; w[42][176] = 5'b10000; w[42][177] = 5'b00000; w[42][178] = 5'b01111; w[42][179] = 5'b01111; w[42][180] = 5'b01111; w[42][181] = 5'b01111; w[42][182] = 5'b01111; w[42][183] = 5'b01111; w[42][184] = 5'b01111; w[42][185] = 5'b01111; w[42][186] = 5'b01111; w[42][187] = 5'b01111; w[42][188] = 5'b01111; w[42][189] = 5'b01111; w[42][190] = 5'b01111; w[42][191] = 5'b01111; w[42][192] = 5'b01111; w[42][193] = 5'b01111; w[42][194] = 5'b01111; w[42][195] = 5'b01111; w[42][196] = 5'b01111; w[42][197] = 5'b01111; w[42][198] = 5'b01111; w[42][199] = 5'b01111; w[42][200] = 5'b01111; w[42][201] = 5'b01111; w[42][202] = 5'b01111; w[42][203] = 5'b01111; w[42][204] = 5'b01111; w[42][205] = 5'b01111; w[42][206] = 5'b01111; w[42][207] = 5'b01111; w[42][208] = 5'b01111; w[42][209] = 5'b01111; 
w[43][0] = 5'b01111; w[43][1] = 5'b01111; w[43][2] = 5'b01111; w[43][3] = 5'b01111; w[43][4] = 5'b01111; w[43][5] = 5'b01111; w[43][6] = 5'b01111; w[43][7] = 5'b01111; w[43][8] = 5'b01111; w[43][9] = 5'b01111; w[43][10] = 5'b01111; w[43][11] = 5'b01111; w[43][12] = 5'b01111; w[43][13] = 5'b01111; w[43][14] = 5'b01111; w[43][15] = 5'b01111; w[43][16] = 5'b01111; w[43][17] = 5'b01111; w[43][18] = 5'b01111; w[43][19] = 5'b01111; w[43][20] = 5'b01111; w[43][21] = 5'b01111; w[43][22] = 5'b01111; w[43][23] = 5'b01111; w[43][24] = 5'b01111; w[43][25] = 5'b01111; w[43][26] = 5'b01111; w[43][27] = 5'b01111; w[43][28] = 5'b01111; w[43][29] = 5'b01111; w[43][30] = 5'b01111; w[43][31] = 5'b00000; w[43][32] = 5'b10000; w[43][33] = 5'b10000; w[43][34] = 5'b10000; w[43][35] = 5'b10000; w[43][36] = 5'b10000; w[43][37] = 5'b10000; w[43][38] = 5'b00000; w[43][39] = 5'b01111; w[43][40] = 5'b01111; w[43][41] = 5'b01111; w[43][42] = 5'b01111; w[43][43] = 5'b00000; w[43][44] = 5'b01111; w[43][45] = 5'b10000; w[43][46] = 5'b10000; w[43][47] = 5'b10000; w[43][48] = 5'b10000; w[43][49] = 5'b10000; w[43][50] = 5'b10000; w[43][51] = 5'b10000; w[43][52] = 5'b10000; w[43][53] = 5'b01111; w[43][54] = 5'b01111; w[43][55] = 5'b01111; w[43][56] = 5'b01111; w[43][57] = 5'b01111; w[43][58] = 5'b01111; w[43][59] = 5'b00000; w[43][60] = 5'b00000; w[43][61] = 5'b01111; w[43][62] = 5'b10000; w[43][63] = 5'b00000; w[43][64] = 5'b01111; w[43][65] = 5'b00000; w[43][66] = 5'b00000; w[43][67] = 5'b01111; w[43][68] = 5'b01111; w[43][69] = 5'b01111; w[43][70] = 5'b01111; w[43][71] = 5'b01111; w[43][72] = 5'b01111; w[43][73] = 5'b00000; w[43][74] = 5'b01111; w[43][75] = 5'b01111; w[43][76] = 5'b10000; w[43][77] = 5'b00000; w[43][78] = 5'b01111; w[43][79] = 5'b01111; w[43][80] = 5'b00000; w[43][81] = 5'b01111; w[43][82] = 5'b01111; w[43][83] = 5'b01111; w[43][84] = 5'b01111; w[43][85] = 5'b01111; w[43][86] = 5'b01111; w[43][87] = 5'b00000; w[43][88] = 5'b01111; w[43][89] = 5'b01111; w[43][90] = 5'b10000; w[43][91] = 5'b10000; w[43][92] = 5'b01111; w[43][93] = 5'b01111; w[43][94] = 5'b01111; w[43][95] = 5'b01111; w[43][96] = 5'b01111; w[43][97] = 5'b01111; w[43][98] = 5'b01111; w[43][99] = 5'b01111; w[43][100] = 5'b01111; w[43][101] = 5'b00000; w[43][102] = 5'b01111; w[43][103] = 5'b01111; w[43][104] = 5'b10000; w[43][105] = 5'b10000; w[43][106] = 5'b01111; w[43][107] = 5'b00000; w[43][108] = 5'b00000; w[43][109] = 5'b01111; w[43][110] = 5'b01111; w[43][111] = 5'b01111; w[43][112] = 5'b01111; w[43][113] = 5'b01111; w[43][114] = 5'b01111; w[43][115] = 5'b00000; w[43][116] = 5'b01111; w[43][117] = 5'b01111; w[43][118] = 5'b10000; w[43][119] = 5'b10000; w[43][120] = 5'b00000; w[43][121] = 5'b00000; w[43][122] = 5'b00000; w[43][123] = 5'b01111; w[43][124] = 5'b01111; w[43][125] = 5'b01111; w[43][126] = 5'b01111; w[43][127] = 5'b01111; w[43][128] = 5'b01111; w[43][129] = 5'b00000; w[43][130] = 5'b01111; w[43][131] = 5'b01111; w[43][132] = 5'b00000; w[43][133] = 5'b10000; w[43][134] = 5'b01111; w[43][135] = 5'b01111; w[43][136] = 5'b00000; w[43][137] = 5'b01111; w[43][138] = 5'b01111; w[43][139] = 5'b01111; w[43][140] = 5'b01111; w[43][141] = 5'b01111; w[43][142] = 5'b01111; w[43][143] = 5'b00000; w[43][144] = 5'b00000; w[43][145] = 5'b01111; w[43][146] = 5'b00000; w[43][147] = 5'b10000; w[43][148] = 5'b01111; w[43][149] = 5'b00000; w[43][150] = 5'b00000; w[43][151] = 5'b01111; w[43][152] = 5'b01111; w[43][153] = 5'b01111; w[43][154] = 5'b01111; w[43][155] = 5'b01111; w[43][156] = 5'b01111; w[43][157] = 5'b00000; w[43][158] = 5'b00000; w[43][159] = 5'b00000; w[43][160] = 5'b10000; w[43][161] = 5'b10000; w[43][162] = 5'b10000; w[43][163] = 5'b00000; w[43][164] = 5'b00000; w[43][165] = 5'b01111; w[43][166] = 5'b01111; w[43][167] = 5'b01111; w[43][168] = 5'b01111; w[43][169] = 5'b01111; w[43][170] = 5'b01111; w[43][171] = 5'b01111; w[43][172] = 5'b00000; w[43][173] = 5'b00000; w[43][174] = 5'b10000; w[43][175] = 5'b10000; w[43][176] = 5'b10000; w[43][177] = 5'b00000; w[43][178] = 5'b01111; w[43][179] = 5'b01111; w[43][180] = 5'b01111; w[43][181] = 5'b01111; w[43][182] = 5'b01111; w[43][183] = 5'b01111; w[43][184] = 5'b01111; w[43][185] = 5'b01111; w[43][186] = 5'b01111; w[43][187] = 5'b01111; w[43][188] = 5'b01111; w[43][189] = 5'b01111; w[43][190] = 5'b01111; w[43][191] = 5'b01111; w[43][192] = 5'b01111; w[43][193] = 5'b01111; w[43][194] = 5'b01111; w[43][195] = 5'b01111; w[43][196] = 5'b01111; w[43][197] = 5'b01111; w[43][198] = 5'b01111; w[43][199] = 5'b01111; w[43][200] = 5'b01111; w[43][201] = 5'b01111; w[43][202] = 5'b01111; w[43][203] = 5'b01111; w[43][204] = 5'b01111; w[43][205] = 5'b01111; w[43][206] = 5'b01111; w[43][207] = 5'b01111; w[43][208] = 5'b01111; w[43][209] = 5'b01111; 
w[44][0] = 5'b01111; w[44][1] = 5'b01111; w[44][2] = 5'b01111; w[44][3] = 5'b01111; w[44][4] = 5'b01111; w[44][5] = 5'b01111; w[44][6] = 5'b01111; w[44][7] = 5'b01111; w[44][8] = 5'b01111; w[44][9] = 5'b01111; w[44][10] = 5'b01111; w[44][11] = 5'b01111; w[44][12] = 5'b01111; w[44][13] = 5'b01111; w[44][14] = 5'b01111; w[44][15] = 5'b01111; w[44][16] = 5'b01111; w[44][17] = 5'b01111; w[44][18] = 5'b01111; w[44][19] = 5'b01111; w[44][20] = 5'b01111; w[44][21] = 5'b01111; w[44][22] = 5'b01111; w[44][23] = 5'b01111; w[44][24] = 5'b01111; w[44][25] = 5'b01111; w[44][26] = 5'b01111; w[44][27] = 5'b01111; w[44][28] = 5'b01111; w[44][29] = 5'b01111; w[44][30] = 5'b01111; w[44][31] = 5'b01111; w[44][32] = 5'b00000; w[44][33] = 5'b10000; w[44][34] = 5'b00000; w[44][35] = 5'b00000; w[44][36] = 5'b00000; w[44][37] = 5'b00000; w[44][38] = 5'b01111; w[44][39] = 5'b01111; w[44][40] = 5'b01111; w[44][41] = 5'b01111; w[44][42] = 5'b01111; w[44][43] = 5'b01111; w[44][44] = 5'b00000; w[44][45] = 5'b00000; w[44][46] = 5'b00000; w[44][47] = 5'b10000; w[44][48] = 5'b00000; w[44][49] = 5'b00000; w[44][50] = 5'b00000; w[44][51] = 5'b00000; w[44][52] = 5'b00000; w[44][53] = 5'b01111; w[44][54] = 5'b01111; w[44][55] = 5'b01111; w[44][56] = 5'b01111; w[44][57] = 5'b01111; w[44][58] = 5'b00000; w[44][59] = 5'b10000; w[44][60] = 5'b10000; w[44][61] = 5'b00000; w[44][62] = 5'b00000; w[44][63] = 5'b01111; w[44][64] = 5'b01111; w[44][65] = 5'b10000; w[44][66] = 5'b10000; w[44][67] = 5'b00000; w[44][68] = 5'b01111; w[44][69] = 5'b01111; w[44][70] = 5'b01111; w[44][71] = 5'b01111; w[44][72] = 5'b00000; w[44][73] = 5'b10000; w[44][74] = 5'b00000; w[44][75] = 5'b00000; w[44][76] = 5'b00000; w[44][77] = 5'b01111; w[44][78] = 5'b01111; w[44][79] = 5'b00000; w[44][80] = 5'b10000; w[44][81] = 5'b00000; w[44][82] = 5'b01111; w[44][83] = 5'b01111; w[44][84] = 5'b01111; w[44][85] = 5'b01111; w[44][86] = 5'b00000; w[44][87] = 5'b10000; w[44][88] = 5'b00000; w[44][89] = 5'b00000; w[44][90] = 5'b00000; w[44][91] = 5'b00000; w[44][92] = 5'b01111; w[44][93] = 5'b00000; w[44][94] = 5'b00000; w[44][95] = 5'b01111; w[44][96] = 5'b01111; w[44][97] = 5'b01111; w[44][98] = 5'b01111; w[44][99] = 5'b01111; w[44][100] = 5'b00000; w[44][101] = 5'b10000; w[44][102] = 5'b00000; w[44][103] = 5'b01111; w[44][104] = 5'b00000; w[44][105] = 5'b00000; w[44][106] = 5'b00000; w[44][107] = 5'b10000; w[44][108] = 5'b10000; w[44][109] = 5'b00000; w[44][110] = 5'b01111; w[44][111] = 5'b01111; w[44][112] = 5'b01111; w[44][113] = 5'b01111; w[44][114] = 5'b00000; w[44][115] = 5'b10000; w[44][116] = 5'b00000; w[44][117] = 5'b01111; w[44][118] = 5'b00000; w[44][119] = 5'b00000; w[44][120] = 5'b10000; w[44][121] = 5'b10000; w[44][122] = 5'b10000; w[44][123] = 5'b00000; w[44][124] = 5'b01111; w[44][125] = 5'b01111; w[44][126] = 5'b01111; w[44][127] = 5'b01111; w[44][128] = 5'b00000; w[44][129] = 5'b10000; w[44][130] = 5'b00000; w[44][131] = 5'b01111; w[44][132] = 5'b01111; w[44][133] = 5'b00000; w[44][134] = 5'b00000; w[44][135] = 5'b00000; w[44][136] = 5'b10000; w[44][137] = 5'b00000; w[44][138] = 5'b01111; w[44][139] = 5'b01111; w[44][140] = 5'b01111; w[44][141] = 5'b01111; w[44][142] = 5'b00000; w[44][143] = 5'b10000; w[44][144] = 5'b10000; w[44][145] = 5'b01111; w[44][146] = 5'b01111; w[44][147] = 5'b00000; w[44][148] = 5'b00000; w[44][149] = 5'b10000; w[44][150] = 5'b10000; w[44][151] = 5'b00000; w[44][152] = 5'b01111; w[44][153] = 5'b01111; w[44][154] = 5'b01111; w[44][155] = 5'b01111; w[44][156] = 5'b01111; w[44][157] = 5'b10000; w[44][158] = 5'b10000; w[44][159] = 5'b10000; w[44][160] = 5'b00000; w[44][161] = 5'b00000; w[44][162] = 5'b10000; w[44][163] = 5'b10000; w[44][164] = 5'b10000; w[44][165] = 5'b01111; w[44][166] = 5'b01111; w[44][167] = 5'b01111; w[44][168] = 5'b01111; w[44][169] = 5'b01111; w[44][170] = 5'b01111; w[44][171] = 5'b00000; w[44][172] = 5'b10000; w[44][173] = 5'b10000; w[44][174] = 5'b00000; w[44][175] = 5'b00000; w[44][176] = 5'b10000; w[44][177] = 5'b10000; w[44][178] = 5'b00000; w[44][179] = 5'b01111; w[44][180] = 5'b01111; w[44][181] = 5'b01111; w[44][182] = 5'b01111; w[44][183] = 5'b01111; w[44][184] = 5'b01111; w[44][185] = 5'b01111; w[44][186] = 5'b01111; w[44][187] = 5'b01111; w[44][188] = 5'b01111; w[44][189] = 5'b01111; w[44][190] = 5'b01111; w[44][191] = 5'b01111; w[44][192] = 5'b01111; w[44][193] = 5'b01111; w[44][194] = 5'b01111; w[44][195] = 5'b01111; w[44][196] = 5'b01111; w[44][197] = 5'b01111; w[44][198] = 5'b01111; w[44][199] = 5'b01111; w[44][200] = 5'b01111; w[44][201] = 5'b01111; w[44][202] = 5'b01111; w[44][203] = 5'b01111; w[44][204] = 5'b01111; w[44][205] = 5'b01111; w[44][206] = 5'b01111; w[44][207] = 5'b01111; w[44][208] = 5'b01111; w[44][209] = 5'b01111; 
w[45][0] = 5'b10000; w[45][1] = 5'b10000; w[45][2] = 5'b10000; w[45][3] = 5'b10000; w[45][4] = 5'b10000; w[45][5] = 5'b10000; w[45][6] = 5'b10000; w[45][7] = 5'b10000; w[45][8] = 5'b10000; w[45][9] = 5'b10000; w[45][10] = 5'b10000; w[45][11] = 5'b10000; w[45][12] = 5'b10000; w[45][13] = 5'b10000; w[45][14] = 5'b10000; w[45][15] = 5'b10000; w[45][16] = 5'b10000; w[45][17] = 5'b10000; w[45][18] = 5'b10000; w[45][19] = 5'b10000; w[45][20] = 5'b10000; w[45][21] = 5'b10000; w[45][22] = 5'b10000; w[45][23] = 5'b10000; w[45][24] = 5'b10000; w[45][25] = 5'b10000; w[45][26] = 5'b10000; w[45][27] = 5'b10000; w[45][28] = 5'b10000; w[45][29] = 5'b10000; w[45][30] = 5'b00000; w[45][31] = 5'b01111; w[45][32] = 5'b01111; w[45][33] = 5'b01111; w[45][34] = 5'b00000; w[45][35] = 5'b00000; w[45][36] = 5'b00000; w[45][37] = 5'b01111; w[45][38] = 5'b01111; w[45][39] = 5'b00000; w[45][40] = 5'b10000; w[45][41] = 5'b10000; w[45][42] = 5'b10000; w[45][43] = 5'b10000; w[45][44] = 5'b00000; w[45][45] = 5'b00000; w[45][46] = 5'b01111; w[45][47] = 5'b01111; w[45][48] = 5'b00000; w[45][49] = 5'b00000; w[45][50] = 5'b00000; w[45][51] = 5'b01111; w[45][52] = 5'b01111; w[45][53] = 5'b00000; w[45][54] = 5'b10000; w[45][55] = 5'b10000; w[45][56] = 5'b10000; w[45][57] = 5'b10000; w[45][58] = 5'b00000; w[45][59] = 5'b01111; w[45][60] = 5'b01111; w[45][61] = 5'b00000; w[45][62] = 5'b00000; w[45][63] = 5'b10000; w[45][64] = 5'b10000; w[45][65] = 5'b01111; w[45][66] = 5'b01111; w[45][67] = 5'b00000; w[45][68] = 5'b10000; w[45][69] = 5'b10000; w[45][70] = 5'b10000; w[45][71] = 5'b10000; w[45][72] = 5'b00000; w[45][73] = 5'b01111; w[45][74] = 5'b00000; w[45][75] = 5'b00000; w[45][76] = 5'b00000; w[45][77] = 5'b10000; w[45][78] = 5'b10000; w[45][79] = 5'b00000; w[45][80] = 5'b01111; w[45][81] = 5'b00000; w[45][82] = 5'b10000; w[45][83] = 5'b10000; w[45][84] = 5'b10000; w[45][85] = 5'b10000; w[45][86] = 5'b00000; w[45][87] = 5'b01111; w[45][88] = 5'b00000; w[45][89] = 5'b00000; w[45][90] = 5'b00000; w[45][91] = 5'b00000; w[45][92] = 5'b10000; w[45][93] = 5'b00000; w[45][94] = 5'b00000; w[45][95] = 5'b10000; w[45][96] = 5'b10000; w[45][97] = 5'b10000; w[45][98] = 5'b10000; w[45][99] = 5'b10000; w[45][100] = 5'b00000; w[45][101] = 5'b01111; w[45][102] = 5'b00000; w[45][103] = 5'b10000; w[45][104] = 5'b00000; w[45][105] = 5'b00000; w[45][106] = 5'b00000; w[45][107] = 5'b01111; w[45][108] = 5'b01111; w[45][109] = 5'b00000; w[45][110] = 5'b10000; w[45][111] = 5'b10000; w[45][112] = 5'b10000; w[45][113] = 5'b10000; w[45][114] = 5'b00000; w[45][115] = 5'b01111; w[45][116] = 5'b00000; w[45][117] = 5'b10000; w[45][118] = 5'b00000; w[45][119] = 5'b00000; w[45][120] = 5'b01111; w[45][121] = 5'b01111; w[45][122] = 5'b01111; w[45][123] = 5'b00000; w[45][124] = 5'b10000; w[45][125] = 5'b10000; w[45][126] = 5'b10000; w[45][127] = 5'b10000; w[45][128] = 5'b00000; w[45][129] = 5'b01111; w[45][130] = 5'b00000; w[45][131] = 5'b10000; w[45][132] = 5'b10000; w[45][133] = 5'b00000; w[45][134] = 5'b00000; w[45][135] = 5'b00000; w[45][136] = 5'b01111; w[45][137] = 5'b00000; w[45][138] = 5'b10000; w[45][139] = 5'b10000; w[45][140] = 5'b10000; w[45][141] = 5'b10000; w[45][142] = 5'b00000; w[45][143] = 5'b01111; w[45][144] = 5'b01111; w[45][145] = 5'b10000; w[45][146] = 5'b10000; w[45][147] = 5'b00000; w[45][148] = 5'b00000; w[45][149] = 5'b01111; w[45][150] = 5'b01111; w[45][151] = 5'b00000; w[45][152] = 5'b10000; w[45][153] = 5'b10000; w[45][154] = 5'b10000; w[45][155] = 5'b10000; w[45][156] = 5'b10000; w[45][157] = 5'b01111; w[45][158] = 5'b01111; w[45][159] = 5'b10000; w[45][160] = 5'b00000; w[45][161] = 5'b00000; w[45][162] = 5'b00000; w[45][163] = 5'b01111; w[45][164] = 5'b01111; w[45][165] = 5'b10000; w[45][166] = 5'b10000; w[45][167] = 5'b10000; w[45][168] = 5'b10000; w[45][169] = 5'b10000; w[45][170] = 5'b10000; w[45][171] = 5'b00000; w[45][172] = 5'b01111; w[45][173] = 5'b10000; w[45][174] = 5'b00000; w[45][175] = 5'b00000; w[45][176] = 5'b00000; w[45][177] = 5'b01111; w[45][178] = 5'b00000; w[45][179] = 5'b10000; w[45][180] = 5'b10000; w[45][181] = 5'b10000; w[45][182] = 5'b10000; w[45][183] = 5'b10000; w[45][184] = 5'b10000; w[45][185] = 5'b10000; w[45][186] = 5'b10000; w[45][187] = 5'b10000; w[45][188] = 5'b10000; w[45][189] = 5'b10000; w[45][190] = 5'b10000; w[45][191] = 5'b10000; w[45][192] = 5'b10000; w[45][193] = 5'b10000; w[45][194] = 5'b10000; w[45][195] = 5'b10000; w[45][196] = 5'b10000; w[45][197] = 5'b10000; w[45][198] = 5'b10000; w[45][199] = 5'b10000; w[45][200] = 5'b10000; w[45][201] = 5'b10000; w[45][202] = 5'b10000; w[45][203] = 5'b10000; w[45][204] = 5'b10000; w[45][205] = 5'b10000; w[45][206] = 5'b10000; w[45][207] = 5'b10000; w[45][208] = 5'b10000; w[45][209] = 5'b10000; 
w[46][0] = 5'b10000; w[46][1] = 5'b10000; w[46][2] = 5'b10000; w[46][3] = 5'b10000; w[46][4] = 5'b10000; w[46][5] = 5'b10000; w[46][6] = 5'b10000; w[46][7] = 5'b10000; w[46][8] = 5'b10000; w[46][9] = 5'b10000; w[46][10] = 5'b10000; w[46][11] = 5'b10000; w[46][12] = 5'b10000; w[46][13] = 5'b10000; w[46][14] = 5'b10000; w[46][15] = 5'b10000; w[46][16] = 5'b10000; w[46][17] = 5'b10000; w[46][18] = 5'b10000; w[46][19] = 5'b10000; w[46][20] = 5'b10000; w[46][21] = 5'b10000; w[46][22] = 5'b10000; w[46][23] = 5'b10000; w[46][24] = 5'b10000; w[46][25] = 5'b10000; w[46][26] = 5'b10000; w[46][27] = 5'b10000; w[46][28] = 5'b10000; w[46][29] = 5'b10000; w[46][30] = 5'b00000; w[46][31] = 5'b01111; w[46][32] = 5'b01111; w[46][33] = 5'b01111; w[46][34] = 5'b00000; w[46][35] = 5'b00000; w[46][36] = 5'b00000; w[46][37] = 5'b01111; w[46][38] = 5'b01111; w[46][39] = 5'b00000; w[46][40] = 5'b10000; w[46][41] = 5'b10000; w[46][42] = 5'b10000; w[46][43] = 5'b10000; w[46][44] = 5'b00000; w[46][45] = 5'b01111; w[46][46] = 5'b00000; w[46][47] = 5'b01111; w[46][48] = 5'b00000; w[46][49] = 5'b00000; w[46][50] = 5'b00000; w[46][51] = 5'b01111; w[46][52] = 5'b01111; w[46][53] = 5'b00000; w[46][54] = 5'b10000; w[46][55] = 5'b10000; w[46][56] = 5'b10000; w[46][57] = 5'b10000; w[46][58] = 5'b00000; w[46][59] = 5'b01111; w[46][60] = 5'b01111; w[46][61] = 5'b00000; w[46][62] = 5'b00000; w[46][63] = 5'b10000; w[46][64] = 5'b10000; w[46][65] = 5'b01111; w[46][66] = 5'b01111; w[46][67] = 5'b00000; w[46][68] = 5'b10000; w[46][69] = 5'b10000; w[46][70] = 5'b10000; w[46][71] = 5'b10000; w[46][72] = 5'b00000; w[46][73] = 5'b01111; w[46][74] = 5'b00000; w[46][75] = 5'b00000; w[46][76] = 5'b00000; w[46][77] = 5'b10000; w[46][78] = 5'b10000; w[46][79] = 5'b00000; w[46][80] = 5'b01111; w[46][81] = 5'b00000; w[46][82] = 5'b10000; w[46][83] = 5'b10000; w[46][84] = 5'b10000; w[46][85] = 5'b10000; w[46][86] = 5'b00000; w[46][87] = 5'b01111; w[46][88] = 5'b00000; w[46][89] = 5'b00000; w[46][90] = 5'b00000; w[46][91] = 5'b00000; w[46][92] = 5'b10000; w[46][93] = 5'b00000; w[46][94] = 5'b00000; w[46][95] = 5'b10000; w[46][96] = 5'b10000; w[46][97] = 5'b10000; w[46][98] = 5'b10000; w[46][99] = 5'b10000; w[46][100] = 5'b00000; w[46][101] = 5'b01111; w[46][102] = 5'b00000; w[46][103] = 5'b10000; w[46][104] = 5'b00000; w[46][105] = 5'b00000; w[46][106] = 5'b00000; w[46][107] = 5'b01111; w[46][108] = 5'b01111; w[46][109] = 5'b00000; w[46][110] = 5'b10000; w[46][111] = 5'b10000; w[46][112] = 5'b10000; w[46][113] = 5'b10000; w[46][114] = 5'b00000; w[46][115] = 5'b01111; w[46][116] = 5'b00000; w[46][117] = 5'b10000; w[46][118] = 5'b00000; w[46][119] = 5'b00000; w[46][120] = 5'b01111; w[46][121] = 5'b01111; w[46][122] = 5'b01111; w[46][123] = 5'b00000; w[46][124] = 5'b10000; w[46][125] = 5'b10000; w[46][126] = 5'b10000; w[46][127] = 5'b10000; w[46][128] = 5'b00000; w[46][129] = 5'b01111; w[46][130] = 5'b00000; w[46][131] = 5'b10000; w[46][132] = 5'b10000; w[46][133] = 5'b00000; w[46][134] = 5'b00000; w[46][135] = 5'b00000; w[46][136] = 5'b01111; w[46][137] = 5'b00000; w[46][138] = 5'b10000; w[46][139] = 5'b10000; w[46][140] = 5'b10000; w[46][141] = 5'b10000; w[46][142] = 5'b00000; w[46][143] = 5'b01111; w[46][144] = 5'b01111; w[46][145] = 5'b10000; w[46][146] = 5'b10000; w[46][147] = 5'b00000; w[46][148] = 5'b00000; w[46][149] = 5'b01111; w[46][150] = 5'b01111; w[46][151] = 5'b00000; w[46][152] = 5'b10000; w[46][153] = 5'b10000; w[46][154] = 5'b10000; w[46][155] = 5'b10000; w[46][156] = 5'b10000; w[46][157] = 5'b01111; w[46][158] = 5'b01111; w[46][159] = 5'b10000; w[46][160] = 5'b00000; w[46][161] = 5'b00000; w[46][162] = 5'b00000; w[46][163] = 5'b01111; w[46][164] = 5'b01111; w[46][165] = 5'b10000; w[46][166] = 5'b10000; w[46][167] = 5'b10000; w[46][168] = 5'b10000; w[46][169] = 5'b10000; w[46][170] = 5'b10000; w[46][171] = 5'b00000; w[46][172] = 5'b01111; w[46][173] = 5'b10000; w[46][174] = 5'b00000; w[46][175] = 5'b00000; w[46][176] = 5'b00000; w[46][177] = 5'b01111; w[46][178] = 5'b00000; w[46][179] = 5'b10000; w[46][180] = 5'b10000; w[46][181] = 5'b10000; w[46][182] = 5'b10000; w[46][183] = 5'b10000; w[46][184] = 5'b10000; w[46][185] = 5'b10000; w[46][186] = 5'b10000; w[46][187] = 5'b10000; w[46][188] = 5'b10000; w[46][189] = 5'b10000; w[46][190] = 5'b10000; w[46][191] = 5'b10000; w[46][192] = 5'b10000; w[46][193] = 5'b10000; w[46][194] = 5'b10000; w[46][195] = 5'b10000; w[46][196] = 5'b10000; w[46][197] = 5'b10000; w[46][198] = 5'b10000; w[46][199] = 5'b10000; w[46][200] = 5'b10000; w[46][201] = 5'b10000; w[46][202] = 5'b10000; w[46][203] = 5'b10000; w[46][204] = 5'b10000; w[46][205] = 5'b10000; w[46][206] = 5'b10000; w[46][207] = 5'b10000; w[46][208] = 5'b10000; w[46][209] = 5'b10000; 
w[47][0] = 5'b10000; w[47][1] = 5'b10000; w[47][2] = 5'b10000; w[47][3] = 5'b10000; w[47][4] = 5'b10000; w[47][5] = 5'b10000; w[47][6] = 5'b10000; w[47][7] = 5'b10000; w[47][8] = 5'b10000; w[47][9] = 5'b10000; w[47][10] = 5'b10000; w[47][11] = 5'b10000; w[47][12] = 5'b10000; w[47][13] = 5'b10000; w[47][14] = 5'b10000; w[47][15] = 5'b10000; w[47][16] = 5'b10000; w[47][17] = 5'b10000; w[47][18] = 5'b10000; w[47][19] = 5'b10000; w[47][20] = 5'b10000; w[47][21] = 5'b10000; w[47][22] = 5'b10000; w[47][23] = 5'b10000; w[47][24] = 5'b10000; w[47][25] = 5'b10000; w[47][26] = 5'b10000; w[47][27] = 5'b10000; w[47][28] = 5'b10000; w[47][29] = 5'b10000; w[47][30] = 5'b10000; w[47][31] = 5'b00000; w[47][32] = 5'b01111; w[47][33] = 5'b01111; w[47][34] = 5'b01111; w[47][35] = 5'b01111; w[47][36] = 5'b01111; w[47][37] = 5'b01111; w[47][38] = 5'b00000; w[47][39] = 5'b10000; w[47][40] = 5'b10000; w[47][41] = 5'b10000; w[47][42] = 5'b10000; w[47][43] = 5'b10000; w[47][44] = 5'b10000; w[47][45] = 5'b01111; w[47][46] = 5'b01111; w[47][47] = 5'b00000; w[47][48] = 5'b01111; w[47][49] = 5'b01111; w[47][50] = 5'b01111; w[47][51] = 5'b01111; w[47][52] = 5'b01111; w[47][53] = 5'b10000; w[47][54] = 5'b10000; w[47][55] = 5'b10000; w[47][56] = 5'b10000; w[47][57] = 5'b10000; w[47][58] = 5'b10000; w[47][59] = 5'b00000; w[47][60] = 5'b00000; w[47][61] = 5'b10000; w[47][62] = 5'b01111; w[47][63] = 5'b00000; w[47][64] = 5'b10000; w[47][65] = 5'b00000; w[47][66] = 5'b00000; w[47][67] = 5'b10000; w[47][68] = 5'b10000; w[47][69] = 5'b10000; w[47][70] = 5'b10000; w[47][71] = 5'b10000; w[47][72] = 5'b10000; w[47][73] = 5'b00000; w[47][74] = 5'b10000; w[47][75] = 5'b10000; w[47][76] = 5'b01111; w[47][77] = 5'b00000; w[47][78] = 5'b10000; w[47][79] = 5'b10000; w[47][80] = 5'b00000; w[47][81] = 5'b10000; w[47][82] = 5'b10000; w[47][83] = 5'b10000; w[47][84] = 5'b10000; w[47][85] = 5'b10000; w[47][86] = 5'b10000; w[47][87] = 5'b00000; w[47][88] = 5'b10000; w[47][89] = 5'b10000; w[47][90] = 5'b01111; w[47][91] = 5'b01111; w[47][92] = 5'b10000; w[47][93] = 5'b10000; w[47][94] = 5'b10000; w[47][95] = 5'b10000; w[47][96] = 5'b10000; w[47][97] = 5'b10000; w[47][98] = 5'b10000; w[47][99] = 5'b10000; w[47][100] = 5'b10000; w[47][101] = 5'b00000; w[47][102] = 5'b10000; w[47][103] = 5'b10000; w[47][104] = 5'b01111; w[47][105] = 5'b01111; w[47][106] = 5'b10000; w[47][107] = 5'b00000; w[47][108] = 5'b00000; w[47][109] = 5'b10000; w[47][110] = 5'b10000; w[47][111] = 5'b10000; w[47][112] = 5'b10000; w[47][113] = 5'b10000; w[47][114] = 5'b10000; w[47][115] = 5'b00000; w[47][116] = 5'b10000; w[47][117] = 5'b10000; w[47][118] = 5'b01111; w[47][119] = 5'b01111; w[47][120] = 5'b00000; w[47][121] = 5'b00000; w[47][122] = 5'b00000; w[47][123] = 5'b10000; w[47][124] = 5'b10000; w[47][125] = 5'b10000; w[47][126] = 5'b10000; w[47][127] = 5'b10000; w[47][128] = 5'b10000; w[47][129] = 5'b00000; w[47][130] = 5'b10000; w[47][131] = 5'b10000; w[47][132] = 5'b00000; w[47][133] = 5'b01111; w[47][134] = 5'b10000; w[47][135] = 5'b10000; w[47][136] = 5'b00000; w[47][137] = 5'b10000; w[47][138] = 5'b10000; w[47][139] = 5'b10000; w[47][140] = 5'b10000; w[47][141] = 5'b10000; w[47][142] = 5'b10000; w[47][143] = 5'b00000; w[47][144] = 5'b00000; w[47][145] = 5'b10000; w[47][146] = 5'b00000; w[47][147] = 5'b01111; w[47][148] = 5'b10000; w[47][149] = 5'b00000; w[47][150] = 5'b00000; w[47][151] = 5'b10000; w[47][152] = 5'b10000; w[47][153] = 5'b10000; w[47][154] = 5'b10000; w[47][155] = 5'b10000; w[47][156] = 5'b10000; w[47][157] = 5'b00000; w[47][158] = 5'b00000; w[47][159] = 5'b00000; w[47][160] = 5'b01111; w[47][161] = 5'b01111; w[47][162] = 5'b01111; w[47][163] = 5'b00000; w[47][164] = 5'b00000; w[47][165] = 5'b10000; w[47][166] = 5'b10000; w[47][167] = 5'b10000; w[47][168] = 5'b10000; w[47][169] = 5'b10000; w[47][170] = 5'b10000; w[47][171] = 5'b10000; w[47][172] = 5'b00000; w[47][173] = 5'b00000; w[47][174] = 5'b01111; w[47][175] = 5'b01111; w[47][176] = 5'b01111; w[47][177] = 5'b00000; w[47][178] = 5'b10000; w[47][179] = 5'b10000; w[47][180] = 5'b10000; w[47][181] = 5'b10000; w[47][182] = 5'b10000; w[47][183] = 5'b10000; w[47][184] = 5'b10000; w[47][185] = 5'b10000; w[47][186] = 5'b10000; w[47][187] = 5'b10000; w[47][188] = 5'b10000; w[47][189] = 5'b10000; w[47][190] = 5'b10000; w[47][191] = 5'b10000; w[47][192] = 5'b10000; w[47][193] = 5'b10000; w[47][194] = 5'b10000; w[47][195] = 5'b10000; w[47][196] = 5'b10000; w[47][197] = 5'b10000; w[47][198] = 5'b10000; w[47][199] = 5'b10000; w[47][200] = 5'b10000; w[47][201] = 5'b10000; w[47][202] = 5'b10000; w[47][203] = 5'b10000; w[47][204] = 5'b10000; w[47][205] = 5'b10000; w[47][206] = 5'b10000; w[47][207] = 5'b10000; w[47][208] = 5'b10000; w[47][209] = 5'b10000; 
w[48][0] = 5'b10000; w[48][1] = 5'b10000; w[48][2] = 5'b10000; w[48][3] = 5'b10000; w[48][4] = 5'b10000; w[48][5] = 5'b10000; w[48][6] = 5'b10000; w[48][7] = 5'b10000; w[48][8] = 5'b10000; w[48][9] = 5'b10000; w[48][10] = 5'b10000; w[48][11] = 5'b10000; w[48][12] = 5'b10000; w[48][13] = 5'b10000; w[48][14] = 5'b10000; w[48][15] = 5'b10000; w[48][16] = 5'b10000; w[48][17] = 5'b10000; w[48][18] = 5'b10000; w[48][19] = 5'b10000; w[48][20] = 5'b10000; w[48][21] = 5'b10000; w[48][22] = 5'b10000; w[48][23] = 5'b10000; w[48][24] = 5'b10000; w[48][25] = 5'b10000; w[48][26] = 5'b10000; w[48][27] = 5'b10000; w[48][28] = 5'b10000; w[48][29] = 5'b10000; w[48][30] = 5'b00000; w[48][31] = 5'b10000; w[48][32] = 5'b00000; w[48][33] = 5'b01111; w[48][34] = 5'b01111; w[48][35] = 5'b01111; w[48][36] = 5'b01111; w[48][37] = 5'b00000; w[48][38] = 5'b10000; w[48][39] = 5'b00000; w[48][40] = 5'b10000; w[48][41] = 5'b10000; w[48][42] = 5'b10000; w[48][43] = 5'b10000; w[48][44] = 5'b00000; w[48][45] = 5'b00000; w[48][46] = 5'b00000; w[48][47] = 5'b01111; w[48][48] = 5'b00000; w[48][49] = 5'b01111; w[48][50] = 5'b01111; w[48][51] = 5'b00000; w[48][52] = 5'b00000; w[48][53] = 5'b00000; w[48][54] = 5'b10000; w[48][55] = 5'b10000; w[48][56] = 5'b10000; w[48][57] = 5'b10000; w[48][58] = 5'b00000; w[48][59] = 5'b10000; w[48][60] = 5'b10000; w[48][61] = 5'b10000; w[48][62] = 5'b00000; w[48][63] = 5'b01111; w[48][64] = 5'b10000; w[48][65] = 5'b10000; w[48][66] = 5'b10000; w[48][67] = 5'b00000; w[48][68] = 5'b10000; w[48][69] = 5'b10000; w[48][70] = 5'b10000; w[48][71] = 5'b10000; w[48][72] = 5'b00000; w[48][73] = 5'b10000; w[48][74] = 5'b10000; w[48][75] = 5'b10000; w[48][76] = 5'b00000; w[48][77] = 5'b01111; w[48][78] = 5'b10000; w[48][79] = 5'b10000; w[48][80] = 5'b10000; w[48][81] = 5'b00000; w[48][82] = 5'b10000; w[48][83] = 5'b10000; w[48][84] = 5'b10000; w[48][85] = 5'b10000; w[48][86] = 5'b00000; w[48][87] = 5'b10000; w[48][88] = 5'b10000; w[48][89] = 5'b10000; w[48][90] = 5'b00000; w[48][91] = 5'b00000; w[48][92] = 5'b10000; w[48][93] = 5'b10000; w[48][94] = 5'b10000; w[48][95] = 5'b10000; w[48][96] = 5'b10000; w[48][97] = 5'b10000; w[48][98] = 5'b10000; w[48][99] = 5'b10000; w[48][100] = 5'b00000; w[48][101] = 5'b10000; w[48][102] = 5'b10000; w[48][103] = 5'b10000; w[48][104] = 5'b00000; w[48][105] = 5'b00000; w[48][106] = 5'b00000; w[48][107] = 5'b10000; w[48][108] = 5'b10000; w[48][109] = 5'b00000; w[48][110] = 5'b10000; w[48][111] = 5'b10000; w[48][112] = 5'b10000; w[48][113] = 5'b10000; w[48][114] = 5'b00000; w[48][115] = 5'b10000; w[48][116] = 5'b10000; w[48][117] = 5'b10000; w[48][118] = 5'b00000; w[48][119] = 5'b00000; w[48][120] = 5'b10000; w[48][121] = 5'b10000; w[48][122] = 5'b10000; w[48][123] = 5'b00000; w[48][124] = 5'b10000; w[48][125] = 5'b10000; w[48][126] = 5'b10000; w[48][127] = 5'b10000; w[48][128] = 5'b00000; w[48][129] = 5'b10000; w[48][130] = 5'b10000; w[48][131] = 5'b10000; w[48][132] = 5'b01111; w[48][133] = 5'b00000; w[48][134] = 5'b10000; w[48][135] = 5'b10000; w[48][136] = 5'b10000; w[48][137] = 5'b00000; w[48][138] = 5'b10000; w[48][139] = 5'b10000; w[48][140] = 5'b10000; w[48][141] = 5'b10000; w[48][142] = 5'b00000; w[48][143] = 5'b10000; w[48][144] = 5'b10000; w[48][145] = 5'b10000; w[48][146] = 5'b01111; w[48][147] = 5'b00000; w[48][148] = 5'b10000; w[48][149] = 5'b10000; w[48][150] = 5'b10000; w[48][151] = 5'b00000; w[48][152] = 5'b10000; w[48][153] = 5'b10000; w[48][154] = 5'b10000; w[48][155] = 5'b10000; w[48][156] = 5'b10000; w[48][157] = 5'b10000; w[48][158] = 5'b10000; w[48][159] = 5'b01111; w[48][160] = 5'b01111; w[48][161] = 5'b01111; w[48][162] = 5'b00000; w[48][163] = 5'b10000; w[48][164] = 5'b10000; w[48][165] = 5'b10000; w[48][166] = 5'b10000; w[48][167] = 5'b10000; w[48][168] = 5'b10000; w[48][169] = 5'b10000; w[48][170] = 5'b10000; w[48][171] = 5'b10000; w[48][172] = 5'b10000; w[48][173] = 5'b01111; w[48][174] = 5'b01111; w[48][175] = 5'b01111; w[48][176] = 5'b00000; w[48][177] = 5'b10000; w[48][178] = 5'b10000; w[48][179] = 5'b10000; w[48][180] = 5'b10000; w[48][181] = 5'b10000; w[48][182] = 5'b10000; w[48][183] = 5'b10000; w[48][184] = 5'b10000; w[48][185] = 5'b10000; w[48][186] = 5'b10000; w[48][187] = 5'b10000; w[48][188] = 5'b10000; w[48][189] = 5'b10000; w[48][190] = 5'b10000; w[48][191] = 5'b10000; w[48][192] = 5'b10000; w[48][193] = 5'b10000; w[48][194] = 5'b10000; w[48][195] = 5'b10000; w[48][196] = 5'b10000; w[48][197] = 5'b10000; w[48][198] = 5'b10000; w[48][199] = 5'b10000; w[48][200] = 5'b10000; w[48][201] = 5'b10000; w[48][202] = 5'b10000; w[48][203] = 5'b10000; w[48][204] = 5'b10000; w[48][205] = 5'b10000; w[48][206] = 5'b10000; w[48][207] = 5'b10000; w[48][208] = 5'b10000; w[48][209] = 5'b10000; 
w[49][0] = 5'b10000; w[49][1] = 5'b10000; w[49][2] = 5'b10000; w[49][3] = 5'b10000; w[49][4] = 5'b10000; w[49][5] = 5'b10000; w[49][6] = 5'b10000; w[49][7] = 5'b10000; w[49][8] = 5'b10000; w[49][9] = 5'b10000; w[49][10] = 5'b10000; w[49][11] = 5'b10000; w[49][12] = 5'b10000; w[49][13] = 5'b10000; w[49][14] = 5'b10000; w[49][15] = 5'b10000; w[49][16] = 5'b10000; w[49][17] = 5'b10000; w[49][18] = 5'b10000; w[49][19] = 5'b10000; w[49][20] = 5'b10000; w[49][21] = 5'b10000; w[49][22] = 5'b10000; w[49][23] = 5'b10000; w[49][24] = 5'b10000; w[49][25] = 5'b10000; w[49][26] = 5'b10000; w[49][27] = 5'b10000; w[49][28] = 5'b10000; w[49][29] = 5'b10000; w[49][30] = 5'b00000; w[49][31] = 5'b10000; w[49][32] = 5'b00000; w[49][33] = 5'b01111; w[49][34] = 5'b01111; w[49][35] = 5'b01111; w[49][36] = 5'b01111; w[49][37] = 5'b00000; w[49][38] = 5'b10000; w[49][39] = 5'b00000; w[49][40] = 5'b10000; w[49][41] = 5'b10000; w[49][42] = 5'b10000; w[49][43] = 5'b10000; w[49][44] = 5'b00000; w[49][45] = 5'b00000; w[49][46] = 5'b00000; w[49][47] = 5'b01111; w[49][48] = 5'b01111; w[49][49] = 5'b00000; w[49][50] = 5'b01111; w[49][51] = 5'b00000; w[49][52] = 5'b00000; w[49][53] = 5'b00000; w[49][54] = 5'b10000; w[49][55] = 5'b10000; w[49][56] = 5'b10000; w[49][57] = 5'b10000; w[49][58] = 5'b00000; w[49][59] = 5'b10000; w[49][60] = 5'b10000; w[49][61] = 5'b10000; w[49][62] = 5'b00000; w[49][63] = 5'b01111; w[49][64] = 5'b10000; w[49][65] = 5'b10000; w[49][66] = 5'b10000; w[49][67] = 5'b00000; w[49][68] = 5'b10000; w[49][69] = 5'b10000; w[49][70] = 5'b10000; w[49][71] = 5'b10000; w[49][72] = 5'b00000; w[49][73] = 5'b10000; w[49][74] = 5'b10000; w[49][75] = 5'b10000; w[49][76] = 5'b00000; w[49][77] = 5'b01111; w[49][78] = 5'b10000; w[49][79] = 5'b10000; w[49][80] = 5'b10000; w[49][81] = 5'b00000; w[49][82] = 5'b10000; w[49][83] = 5'b10000; w[49][84] = 5'b10000; w[49][85] = 5'b10000; w[49][86] = 5'b00000; w[49][87] = 5'b10000; w[49][88] = 5'b10000; w[49][89] = 5'b10000; w[49][90] = 5'b00000; w[49][91] = 5'b00000; w[49][92] = 5'b10000; w[49][93] = 5'b10000; w[49][94] = 5'b10000; w[49][95] = 5'b10000; w[49][96] = 5'b10000; w[49][97] = 5'b10000; w[49][98] = 5'b10000; w[49][99] = 5'b10000; w[49][100] = 5'b00000; w[49][101] = 5'b10000; w[49][102] = 5'b10000; w[49][103] = 5'b10000; w[49][104] = 5'b00000; w[49][105] = 5'b00000; w[49][106] = 5'b00000; w[49][107] = 5'b10000; w[49][108] = 5'b10000; w[49][109] = 5'b00000; w[49][110] = 5'b10000; w[49][111] = 5'b10000; w[49][112] = 5'b10000; w[49][113] = 5'b10000; w[49][114] = 5'b00000; w[49][115] = 5'b10000; w[49][116] = 5'b10000; w[49][117] = 5'b10000; w[49][118] = 5'b00000; w[49][119] = 5'b00000; w[49][120] = 5'b10000; w[49][121] = 5'b10000; w[49][122] = 5'b10000; w[49][123] = 5'b00000; w[49][124] = 5'b10000; w[49][125] = 5'b10000; w[49][126] = 5'b10000; w[49][127] = 5'b10000; w[49][128] = 5'b00000; w[49][129] = 5'b10000; w[49][130] = 5'b10000; w[49][131] = 5'b10000; w[49][132] = 5'b01111; w[49][133] = 5'b00000; w[49][134] = 5'b10000; w[49][135] = 5'b10000; w[49][136] = 5'b10000; w[49][137] = 5'b00000; w[49][138] = 5'b10000; w[49][139] = 5'b10000; w[49][140] = 5'b10000; w[49][141] = 5'b10000; w[49][142] = 5'b00000; w[49][143] = 5'b10000; w[49][144] = 5'b10000; w[49][145] = 5'b10000; w[49][146] = 5'b01111; w[49][147] = 5'b00000; w[49][148] = 5'b10000; w[49][149] = 5'b10000; w[49][150] = 5'b10000; w[49][151] = 5'b00000; w[49][152] = 5'b10000; w[49][153] = 5'b10000; w[49][154] = 5'b10000; w[49][155] = 5'b10000; w[49][156] = 5'b10000; w[49][157] = 5'b10000; w[49][158] = 5'b10000; w[49][159] = 5'b01111; w[49][160] = 5'b01111; w[49][161] = 5'b01111; w[49][162] = 5'b00000; w[49][163] = 5'b10000; w[49][164] = 5'b10000; w[49][165] = 5'b10000; w[49][166] = 5'b10000; w[49][167] = 5'b10000; w[49][168] = 5'b10000; w[49][169] = 5'b10000; w[49][170] = 5'b10000; w[49][171] = 5'b10000; w[49][172] = 5'b10000; w[49][173] = 5'b01111; w[49][174] = 5'b01111; w[49][175] = 5'b01111; w[49][176] = 5'b00000; w[49][177] = 5'b10000; w[49][178] = 5'b10000; w[49][179] = 5'b10000; w[49][180] = 5'b10000; w[49][181] = 5'b10000; w[49][182] = 5'b10000; w[49][183] = 5'b10000; w[49][184] = 5'b10000; w[49][185] = 5'b10000; w[49][186] = 5'b10000; w[49][187] = 5'b10000; w[49][188] = 5'b10000; w[49][189] = 5'b10000; w[49][190] = 5'b10000; w[49][191] = 5'b10000; w[49][192] = 5'b10000; w[49][193] = 5'b10000; w[49][194] = 5'b10000; w[49][195] = 5'b10000; w[49][196] = 5'b10000; w[49][197] = 5'b10000; w[49][198] = 5'b10000; w[49][199] = 5'b10000; w[49][200] = 5'b10000; w[49][201] = 5'b10000; w[49][202] = 5'b10000; w[49][203] = 5'b10000; w[49][204] = 5'b10000; w[49][205] = 5'b10000; w[49][206] = 5'b10000; w[49][207] = 5'b10000; w[49][208] = 5'b10000; w[49][209] = 5'b10000; 
w[50][0] = 5'b10000; w[50][1] = 5'b10000; w[50][2] = 5'b10000; w[50][3] = 5'b10000; w[50][4] = 5'b10000; w[50][5] = 5'b10000; w[50][6] = 5'b10000; w[50][7] = 5'b10000; w[50][8] = 5'b10000; w[50][9] = 5'b10000; w[50][10] = 5'b10000; w[50][11] = 5'b10000; w[50][12] = 5'b10000; w[50][13] = 5'b10000; w[50][14] = 5'b10000; w[50][15] = 5'b10000; w[50][16] = 5'b10000; w[50][17] = 5'b10000; w[50][18] = 5'b10000; w[50][19] = 5'b10000; w[50][20] = 5'b10000; w[50][21] = 5'b10000; w[50][22] = 5'b10000; w[50][23] = 5'b10000; w[50][24] = 5'b10000; w[50][25] = 5'b10000; w[50][26] = 5'b10000; w[50][27] = 5'b10000; w[50][28] = 5'b10000; w[50][29] = 5'b10000; w[50][30] = 5'b00000; w[50][31] = 5'b10000; w[50][32] = 5'b00000; w[50][33] = 5'b01111; w[50][34] = 5'b01111; w[50][35] = 5'b01111; w[50][36] = 5'b01111; w[50][37] = 5'b00000; w[50][38] = 5'b10000; w[50][39] = 5'b00000; w[50][40] = 5'b10000; w[50][41] = 5'b10000; w[50][42] = 5'b10000; w[50][43] = 5'b10000; w[50][44] = 5'b00000; w[50][45] = 5'b00000; w[50][46] = 5'b00000; w[50][47] = 5'b01111; w[50][48] = 5'b01111; w[50][49] = 5'b01111; w[50][50] = 5'b00000; w[50][51] = 5'b00000; w[50][52] = 5'b00000; w[50][53] = 5'b00000; w[50][54] = 5'b10000; w[50][55] = 5'b10000; w[50][56] = 5'b10000; w[50][57] = 5'b10000; w[50][58] = 5'b00000; w[50][59] = 5'b10000; w[50][60] = 5'b10000; w[50][61] = 5'b10000; w[50][62] = 5'b00000; w[50][63] = 5'b01111; w[50][64] = 5'b10000; w[50][65] = 5'b10000; w[50][66] = 5'b10000; w[50][67] = 5'b00000; w[50][68] = 5'b10000; w[50][69] = 5'b10000; w[50][70] = 5'b10000; w[50][71] = 5'b10000; w[50][72] = 5'b00000; w[50][73] = 5'b10000; w[50][74] = 5'b10000; w[50][75] = 5'b10000; w[50][76] = 5'b00000; w[50][77] = 5'b01111; w[50][78] = 5'b10000; w[50][79] = 5'b10000; w[50][80] = 5'b10000; w[50][81] = 5'b00000; w[50][82] = 5'b10000; w[50][83] = 5'b10000; w[50][84] = 5'b10000; w[50][85] = 5'b10000; w[50][86] = 5'b00000; w[50][87] = 5'b10000; w[50][88] = 5'b10000; w[50][89] = 5'b10000; w[50][90] = 5'b00000; w[50][91] = 5'b00000; w[50][92] = 5'b10000; w[50][93] = 5'b10000; w[50][94] = 5'b10000; w[50][95] = 5'b10000; w[50][96] = 5'b10000; w[50][97] = 5'b10000; w[50][98] = 5'b10000; w[50][99] = 5'b10000; w[50][100] = 5'b00000; w[50][101] = 5'b10000; w[50][102] = 5'b10000; w[50][103] = 5'b10000; w[50][104] = 5'b00000; w[50][105] = 5'b00000; w[50][106] = 5'b00000; w[50][107] = 5'b10000; w[50][108] = 5'b10000; w[50][109] = 5'b00000; w[50][110] = 5'b10000; w[50][111] = 5'b10000; w[50][112] = 5'b10000; w[50][113] = 5'b10000; w[50][114] = 5'b00000; w[50][115] = 5'b10000; w[50][116] = 5'b10000; w[50][117] = 5'b10000; w[50][118] = 5'b00000; w[50][119] = 5'b00000; w[50][120] = 5'b10000; w[50][121] = 5'b10000; w[50][122] = 5'b10000; w[50][123] = 5'b00000; w[50][124] = 5'b10000; w[50][125] = 5'b10000; w[50][126] = 5'b10000; w[50][127] = 5'b10000; w[50][128] = 5'b00000; w[50][129] = 5'b10000; w[50][130] = 5'b10000; w[50][131] = 5'b10000; w[50][132] = 5'b01111; w[50][133] = 5'b00000; w[50][134] = 5'b10000; w[50][135] = 5'b10000; w[50][136] = 5'b10000; w[50][137] = 5'b00000; w[50][138] = 5'b10000; w[50][139] = 5'b10000; w[50][140] = 5'b10000; w[50][141] = 5'b10000; w[50][142] = 5'b00000; w[50][143] = 5'b10000; w[50][144] = 5'b10000; w[50][145] = 5'b10000; w[50][146] = 5'b01111; w[50][147] = 5'b00000; w[50][148] = 5'b10000; w[50][149] = 5'b10000; w[50][150] = 5'b10000; w[50][151] = 5'b00000; w[50][152] = 5'b10000; w[50][153] = 5'b10000; w[50][154] = 5'b10000; w[50][155] = 5'b10000; w[50][156] = 5'b10000; w[50][157] = 5'b10000; w[50][158] = 5'b10000; w[50][159] = 5'b01111; w[50][160] = 5'b01111; w[50][161] = 5'b01111; w[50][162] = 5'b00000; w[50][163] = 5'b10000; w[50][164] = 5'b10000; w[50][165] = 5'b10000; w[50][166] = 5'b10000; w[50][167] = 5'b10000; w[50][168] = 5'b10000; w[50][169] = 5'b10000; w[50][170] = 5'b10000; w[50][171] = 5'b10000; w[50][172] = 5'b10000; w[50][173] = 5'b01111; w[50][174] = 5'b01111; w[50][175] = 5'b01111; w[50][176] = 5'b00000; w[50][177] = 5'b10000; w[50][178] = 5'b10000; w[50][179] = 5'b10000; w[50][180] = 5'b10000; w[50][181] = 5'b10000; w[50][182] = 5'b10000; w[50][183] = 5'b10000; w[50][184] = 5'b10000; w[50][185] = 5'b10000; w[50][186] = 5'b10000; w[50][187] = 5'b10000; w[50][188] = 5'b10000; w[50][189] = 5'b10000; w[50][190] = 5'b10000; w[50][191] = 5'b10000; w[50][192] = 5'b10000; w[50][193] = 5'b10000; w[50][194] = 5'b10000; w[50][195] = 5'b10000; w[50][196] = 5'b10000; w[50][197] = 5'b10000; w[50][198] = 5'b10000; w[50][199] = 5'b10000; w[50][200] = 5'b10000; w[50][201] = 5'b10000; w[50][202] = 5'b10000; w[50][203] = 5'b10000; w[50][204] = 5'b10000; w[50][205] = 5'b10000; w[50][206] = 5'b10000; w[50][207] = 5'b10000; w[50][208] = 5'b10000; w[50][209] = 5'b10000; 
w[51][0] = 5'b10000; w[51][1] = 5'b10000; w[51][2] = 5'b10000; w[51][3] = 5'b10000; w[51][4] = 5'b10000; w[51][5] = 5'b10000; w[51][6] = 5'b10000; w[51][7] = 5'b10000; w[51][8] = 5'b10000; w[51][9] = 5'b10000; w[51][10] = 5'b10000; w[51][11] = 5'b10000; w[51][12] = 5'b10000; w[51][13] = 5'b10000; w[51][14] = 5'b10000; w[51][15] = 5'b10000; w[51][16] = 5'b10000; w[51][17] = 5'b10000; w[51][18] = 5'b10000; w[51][19] = 5'b10000; w[51][20] = 5'b10000; w[51][21] = 5'b10000; w[51][22] = 5'b10000; w[51][23] = 5'b10000; w[51][24] = 5'b10000; w[51][25] = 5'b10000; w[51][26] = 5'b10000; w[51][27] = 5'b10000; w[51][28] = 5'b10000; w[51][29] = 5'b10000; w[51][30] = 5'b00000; w[51][31] = 5'b01111; w[51][32] = 5'b01111; w[51][33] = 5'b01111; w[51][34] = 5'b00000; w[51][35] = 5'b00000; w[51][36] = 5'b00000; w[51][37] = 5'b01111; w[51][38] = 5'b01111; w[51][39] = 5'b00000; w[51][40] = 5'b10000; w[51][41] = 5'b10000; w[51][42] = 5'b10000; w[51][43] = 5'b10000; w[51][44] = 5'b00000; w[51][45] = 5'b01111; w[51][46] = 5'b01111; w[51][47] = 5'b01111; w[51][48] = 5'b00000; w[51][49] = 5'b00000; w[51][50] = 5'b00000; w[51][51] = 5'b00000; w[51][52] = 5'b01111; w[51][53] = 5'b00000; w[51][54] = 5'b10000; w[51][55] = 5'b10000; w[51][56] = 5'b10000; w[51][57] = 5'b10000; w[51][58] = 5'b00000; w[51][59] = 5'b01111; w[51][60] = 5'b01111; w[51][61] = 5'b00000; w[51][62] = 5'b00000; w[51][63] = 5'b10000; w[51][64] = 5'b10000; w[51][65] = 5'b01111; w[51][66] = 5'b01111; w[51][67] = 5'b00000; w[51][68] = 5'b10000; w[51][69] = 5'b10000; w[51][70] = 5'b10000; w[51][71] = 5'b10000; w[51][72] = 5'b00000; w[51][73] = 5'b01111; w[51][74] = 5'b00000; w[51][75] = 5'b00000; w[51][76] = 5'b00000; w[51][77] = 5'b10000; w[51][78] = 5'b10000; w[51][79] = 5'b00000; w[51][80] = 5'b01111; w[51][81] = 5'b00000; w[51][82] = 5'b10000; w[51][83] = 5'b10000; w[51][84] = 5'b10000; w[51][85] = 5'b10000; w[51][86] = 5'b00000; w[51][87] = 5'b01111; w[51][88] = 5'b00000; w[51][89] = 5'b00000; w[51][90] = 5'b00000; w[51][91] = 5'b00000; w[51][92] = 5'b10000; w[51][93] = 5'b00000; w[51][94] = 5'b00000; w[51][95] = 5'b10000; w[51][96] = 5'b10000; w[51][97] = 5'b10000; w[51][98] = 5'b10000; w[51][99] = 5'b10000; w[51][100] = 5'b00000; w[51][101] = 5'b01111; w[51][102] = 5'b00000; w[51][103] = 5'b10000; w[51][104] = 5'b00000; w[51][105] = 5'b00000; w[51][106] = 5'b00000; w[51][107] = 5'b01111; w[51][108] = 5'b01111; w[51][109] = 5'b00000; w[51][110] = 5'b10000; w[51][111] = 5'b10000; w[51][112] = 5'b10000; w[51][113] = 5'b10000; w[51][114] = 5'b00000; w[51][115] = 5'b01111; w[51][116] = 5'b00000; w[51][117] = 5'b10000; w[51][118] = 5'b00000; w[51][119] = 5'b00000; w[51][120] = 5'b01111; w[51][121] = 5'b01111; w[51][122] = 5'b01111; w[51][123] = 5'b00000; w[51][124] = 5'b10000; w[51][125] = 5'b10000; w[51][126] = 5'b10000; w[51][127] = 5'b10000; w[51][128] = 5'b00000; w[51][129] = 5'b01111; w[51][130] = 5'b00000; w[51][131] = 5'b10000; w[51][132] = 5'b10000; w[51][133] = 5'b00000; w[51][134] = 5'b00000; w[51][135] = 5'b00000; w[51][136] = 5'b01111; w[51][137] = 5'b00000; w[51][138] = 5'b10000; w[51][139] = 5'b10000; w[51][140] = 5'b10000; w[51][141] = 5'b10000; w[51][142] = 5'b00000; w[51][143] = 5'b01111; w[51][144] = 5'b01111; w[51][145] = 5'b10000; w[51][146] = 5'b10000; w[51][147] = 5'b00000; w[51][148] = 5'b00000; w[51][149] = 5'b01111; w[51][150] = 5'b01111; w[51][151] = 5'b00000; w[51][152] = 5'b10000; w[51][153] = 5'b10000; w[51][154] = 5'b10000; w[51][155] = 5'b10000; w[51][156] = 5'b10000; w[51][157] = 5'b01111; w[51][158] = 5'b01111; w[51][159] = 5'b10000; w[51][160] = 5'b00000; w[51][161] = 5'b00000; w[51][162] = 5'b00000; w[51][163] = 5'b01111; w[51][164] = 5'b01111; w[51][165] = 5'b10000; w[51][166] = 5'b10000; w[51][167] = 5'b10000; w[51][168] = 5'b10000; w[51][169] = 5'b10000; w[51][170] = 5'b10000; w[51][171] = 5'b00000; w[51][172] = 5'b01111; w[51][173] = 5'b10000; w[51][174] = 5'b00000; w[51][175] = 5'b00000; w[51][176] = 5'b00000; w[51][177] = 5'b01111; w[51][178] = 5'b00000; w[51][179] = 5'b10000; w[51][180] = 5'b10000; w[51][181] = 5'b10000; w[51][182] = 5'b10000; w[51][183] = 5'b10000; w[51][184] = 5'b10000; w[51][185] = 5'b10000; w[51][186] = 5'b10000; w[51][187] = 5'b10000; w[51][188] = 5'b10000; w[51][189] = 5'b10000; w[51][190] = 5'b10000; w[51][191] = 5'b10000; w[51][192] = 5'b10000; w[51][193] = 5'b10000; w[51][194] = 5'b10000; w[51][195] = 5'b10000; w[51][196] = 5'b10000; w[51][197] = 5'b10000; w[51][198] = 5'b10000; w[51][199] = 5'b10000; w[51][200] = 5'b10000; w[51][201] = 5'b10000; w[51][202] = 5'b10000; w[51][203] = 5'b10000; w[51][204] = 5'b10000; w[51][205] = 5'b10000; w[51][206] = 5'b10000; w[51][207] = 5'b10000; w[51][208] = 5'b10000; w[51][209] = 5'b10000; 
w[52][0] = 5'b10000; w[52][1] = 5'b10000; w[52][2] = 5'b10000; w[52][3] = 5'b10000; w[52][4] = 5'b10000; w[52][5] = 5'b10000; w[52][6] = 5'b10000; w[52][7] = 5'b10000; w[52][8] = 5'b10000; w[52][9] = 5'b10000; w[52][10] = 5'b10000; w[52][11] = 5'b10000; w[52][12] = 5'b10000; w[52][13] = 5'b10000; w[52][14] = 5'b10000; w[52][15] = 5'b10000; w[52][16] = 5'b10000; w[52][17] = 5'b10000; w[52][18] = 5'b10000; w[52][19] = 5'b10000; w[52][20] = 5'b10000; w[52][21] = 5'b10000; w[52][22] = 5'b10000; w[52][23] = 5'b10000; w[52][24] = 5'b10000; w[52][25] = 5'b10000; w[52][26] = 5'b10000; w[52][27] = 5'b10000; w[52][28] = 5'b10000; w[52][29] = 5'b10000; w[52][30] = 5'b00000; w[52][31] = 5'b01111; w[52][32] = 5'b01111; w[52][33] = 5'b01111; w[52][34] = 5'b00000; w[52][35] = 5'b00000; w[52][36] = 5'b00000; w[52][37] = 5'b01111; w[52][38] = 5'b01111; w[52][39] = 5'b00000; w[52][40] = 5'b10000; w[52][41] = 5'b10000; w[52][42] = 5'b10000; w[52][43] = 5'b10000; w[52][44] = 5'b00000; w[52][45] = 5'b01111; w[52][46] = 5'b01111; w[52][47] = 5'b01111; w[52][48] = 5'b00000; w[52][49] = 5'b00000; w[52][50] = 5'b00000; w[52][51] = 5'b01111; w[52][52] = 5'b00000; w[52][53] = 5'b00000; w[52][54] = 5'b10000; w[52][55] = 5'b10000; w[52][56] = 5'b10000; w[52][57] = 5'b10000; w[52][58] = 5'b00000; w[52][59] = 5'b01111; w[52][60] = 5'b01111; w[52][61] = 5'b00000; w[52][62] = 5'b00000; w[52][63] = 5'b10000; w[52][64] = 5'b10000; w[52][65] = 5'b01111; w[52][66] = 5'b01111; w[52][67] = 5'b00000; w[52][68] = 5'b10000; w[52][69] = 5'b10000; w[52][70] = 5'b10000; w[52][71] = 5'b10000; w[52][72] = 5'b00000; w[52][73] = 5'b01111; w[52][74] = 5'b00000; w[52][75] = 5'b00000; w[52][76] = 5'b00000; w[52][77] = 5'b10000; w[52][78] = 5'b10000; w[52][79] = 5'b00000; w[52][80] = 5'b01111; w[52][81] = 5'b00000; w[52][82] = 5'b10000; w[52][83] = 5'b10000; w[52][84] = 5'b10000; w[52][85] = 5'b10000; w[52][86] = 5'b00000; w[52][87] = 5'b01111; w[52][88] = 5'b00000; w[52][89] = 5'b00000; w[52][90] = 5'b00000; w[52][91] = 5'b00000; w[52][92] = 5'b10000; w[52][93] = 5'b00000; w[52][94] = 5'b00000; w[52][95] = 5'b10000; w[52][96] = 5'b10000; w[52][97] = 5'b10000; w[52][98] = 5'b10000; w[52][99] = 5'b10000; w[52][100] = 5'b00000; w[52][101] = 5'b01111; w[52][102] = 5'b00000; w[52][103] = 5'b10000; w[52][104] = 5'b00000; w[52][105] = 5'b00000; w[52][106] = 5'b00000; w[52][107] = 5'b01111; w[52][108] = 5'b01111; w[52][109] = 5'b00000; w[52][110] = 5'b10000; w[52][111] = 5'b10000; w[52][112] = 5'b10000; w[52][113] = 5'b10000; w[52][114] = 5'b00000; w[52][115] = 5'b01111; w[52][116] = 5'b00000; w[52][117] = 5'b10000; w[52][118] = 5'b00000; w[52][119] = 5'b00000; w[52][120] = 5'b01111; w[52][121] = 5'b01111; w[52][122] = 5'b01111; w[52][123] = 5'b00000; w[52][124] = 5'b10000; w[52][125] = 5'b10000; w[52][126] = 5'b10000; w[52][127] = 5'b10000; w[52][128] = 5'b00000; w[52][129] = 5'b01111; w[52][130] = 5'b00000; w[52][131] = 5'b10000; w[52][132] = 5'b10000; w[52][133] = 5'b00000; w[52][134] = 5'b00000; w[52][135] = 5'b00000; w[52][136] = 5'b01111; w[52][137] = 5'b00000; w[52][138] = 5'b10000; w[52][139] = 5'b10000; w[52][140] = 5'b10000; w[52][141] = 5'b10000; w[52][142] = 5'b00000; w[52][143] = 5'b01111; w[52][144] = 5'b01111; w[52][145] = 5'b10000; w[52][146] = 5'b10000; w[52][147] = 5'b00000; w[52][148] = 5'b00000; w[52][149] = 5'b01111; w[52][150] = 5'b01111; w[52][151] = 5'b00000; w[52][152] = 5'b10000; w[52][153] = 5'b10000; w[52][154] = 5'b10000; w[52][155] = 5'b10000; w[52][156] = 5'b10000; w[52][157] = 5'b01111; w[52][158] = 5'b01111; w[52][159] = 5'b10000; w[52][160] = 5'b00000; w[52][161] = 5'b00000; w[52][162] = 5'b00000; w[52][163] = 5'b01111; w[52][164] = 5'b01111; w[52][165] = 5'b10000; w[52][166] = 5'b10000; w[52][167] = 5'b10000; w[52][168] = 5'b10000; w[52][169] = 5'b10000; w[52][170] = 5'b10000; w[52][171] = 5'b00000; w[52][172] = 5'b01111; w[52][173] = 5'b10000; w[52][174] = 5'b00000; w[52][175] = 5'b00000; w[52][176] = 5'b00000; w[52][177] = 5'b01111; w[52][178] = 5'b00000; w[52][179] = 5'b10000; w[52][180] = 5'b10000; w[52][181] = 5'b10000; w[52][182] = 5'b10000; w[52][183] = 5'b10000; w[52][184] = 5'b10000; w[52][185] = 5'b10000; w[52][186] = 5'b10000; w[52][187] = 5'b10000; w[52][188] = 5'b10000; w[52][189] = 5'b10000; w[52][190] = 5'b10000; w[52][191] = 5'b10000; w[52][192] = 5'b10000; w[52][193] = 5'b10000; w[52][194] = 5'b10000; w[52][195] = 5'b10000; w[52][196] = 5'b10000; w[52][197] = 5'b10000; w[52][198] = 5'b10000; w[52][199] = 5'b10000; w[52][200] = 5'b10000; w[52][201] = 5'b10000; w[52][202] = 5'b10000; w[52][203] = 5'b10000; w[52][204] = 5'b10000; w[52][205] = 5'b10000; w[52][206] = 5'b10000; w[52][207] = 5'b10000; w[52][208] = 5'b10000; w[52][209] = 5'b10000; 
w[53][0] = 5'b01111; w[53][1] = 5'b01111; w[53][2] = 5'b01111; w[53][3] = 5'b01111; w[53][4] = 5'b01111; w[53][5] = 5'b01111; w[53][6] = 5'b01111; w[53][7] = 5'b01111; w[53][8] = 5'b01111; w[53][9] = 5'b01111; w[53][10] = 5'b01111; w[53][11] = 5'b01111; w[53][12] = 5'b01111; w[53][13] = 5'b01111; w[53][14] = 5'b01111; w[53][15] = 5'b01111; w[53][16] = 5'b01111; w[53][17] = 5'b01111; w[53][18] = 5'b01111; w[53][19] = 5'b01111; w[53][20] = 5'b01111; w[53][21] = 5'b01111; w[53][22] = 5'b01111; w[53][23] = 5'b01111; w[53][24] = 5'b01111; w[53][25] = 5'b01111; w[53][26] = 5'b01111; w[53][27] = 5'b01111; w[53][28] = 5'b01111; w[53][29] = 5'b01111; w[53][30] = 5'b01111; w[53][31] = 5'b01111; w[53][32] = 5'b00000; w[53][33] = 5'b10000; w[53][34] = 5'b00000; w[53][35] = 5'b00000; w[53][36] = 5'b00000; w[53][37] = 5'b00000; w[53][38] = 5'b01111; w[53][39] = 5'b01111; w[53][40] = 5'b01111; w[53][41] = 5'b01111; w[53][42] = 5'b01111; w[53][43] = 5'b01111; w[53][44] = 5'b01111; w[53][45] = 5'b00000; w[53][46] = 5'b00000; w[53][47] = 5'b10000; w[53][48] = 5'b00000; w[53][49] = 5'b00000; w[53][50] = 5'b00000; w[53][51] = 5'b00000; w[53][52] = 5'b00000; w[53][53] = 5'b00000; w[53][54] = 5'b01111; w[53][55] = 5'b01111; w[53][56] = 5'b01111; w[53][57] = 5'b01111; w[53][58] = 5'b00000; w[53][59] = 5'b10000; w[53][60] = 5'b10000; w[53][61] = 5'b00000; w[53][62] = 5'b00000; w[53][63] = 5'b01111; w[53][64] = 5'b01111; w[53][65] = 5'b10000; w[53][66] = 5'b10000; w[53][67] = 5'b00000; w[53][68] = 5'b01111; w[53][69] = 5'b01111; w[53][70] = 5'b01111; w[53][71] = 5'b01111; w[53][72] = 5'b00000; w[53][73] = 5'b10000; w[53][74] = 5'b00000; w[53][75] = 5'b00000; w[53][76] = 5'b00000; w[53][77] = 5'b01111; w[53][78] = 5'b01111; w[53][79] = 5'b00000; w[53][80] = 5'b10000; w[53][81] = 5'b00000; w[53][82] = 5'b01111; w[53][83] = 5'b01111; w[53][84] = 5'b01111; w[53][85] = 5'b01111; w[53][86] = 5'b00000; w[53][87] = 5'b10000; w[53][88] = 5'b00000; w[53][89] = 5'b00000; w[53][90] = 5'b00000; w[53][91] = 5'b00000; w[53][92] = 5'b01111; w[53][93] = 5'b00000; w[53][94] = 5'b00000; w[53][95] = 5'b01111; w[53][96] = 5'b01111; w[53][97] = 5'b01111; w[53][98] = 5'b01111; w[53][99] = 5'b01111; w[53][100] = 5'b00000; w[53][101] = 5'b10000; w[53][102] = 5'b00000; w[53][103] = 5'b01111; w[53][104] = 5'b00000; w[53][105] = 5'b00000; w[53][106] = 5'b00000; w[53][107] = 5'b10000; w[53][108] = 5'b10000; w[53][109] = 5'b00000; w[53][110] = 5'b01111; w[53][111] = 5'b01111; w[53][112] = 5'b01111; w[53][113] = 5'b01111; w[53][114] = 5'b00000; w[53][115] = 5'b10000; w[53][116] = 5'b00000; w[53][117] = 5'b01111; w[53][118] = 5'b00000; w[53][119] = 5'b00000; w[53][120] = 5'b10000; w[53][121] = 5'b10000; w[53][122] = 5'b10000; w[53][123] = 5'b00000; w[53][124] = 5'b01111; w[53][125] = 5'b01111; w[53][126] = 5'b01111; w[53][127] = 5'b01111; w[53][128] = 5'b00000; w[53][129] = 5'b10000; w[53][130] = 5'b00000; w[53][131] = 5'b01111; w[53][132] = 5'b01111; w[53][133] = 5'b00000; w[53][134] = 5'b00000; w[53][135] = 5'b00000; w[53][136] = 5'b10000; w[53][137] = 5'b00000; w[53][138] = 5'b01111; w[53][139] = 5'b01111; w[53][140] = 5'b01111; w[53][141] = 5'b01111; w[53][142] = 5'b00000; w[53][143] = 5'b10000; w[53][144] = 5'b10000; w[53][145] = 5'b01111; w[53][146] = 5'b01111; w[53][147] = 5'b00000; w[53][148] = 5'b00000; w[53][149] = 5'b10000; w[53][150] = 5'b10000; w[53][151] = 5'b00000; w[53][152] = 5'b01111; w[53][153] = 5'b01111; w[53][154] = 5'b01111; w[53][155] = 5'b01111; w[53][156] = 5'b01111; w[53][157] = 5'b10000; w[53][158] = 5'b10000; w[53][159] = 5'b10000; w[53][160] = 5'b00000; w[53][161] = 5'b00000; w[53][162] = 5'b10000; w[53][163] = 5'b10000; w[53][164] = 5'b10000; w[53][165] = 5'b01111; w[53][166] = 5'b01111; w[53][167] = 5'b01111; w[53][168] = 5'b01111; w[53][169] = 5'b01111; w[53][170] = 5'b01111; w[53][171] = 5'b00000; w[53][172] = 5'b10000; w[53][173] = 5'b10000; w[53][174] = 5'b00000; w[53][175] = 5'b00000; w[53][176] = 5'b10000; w[53][177] = 5'b10000; w[53][178] = 5'b00000; w[53][179] = 5'b01111; w[53][180] = 5'b01111; w[53][181] = 5'b01111; w[53][182] = 5'b01111; w[53][183] = 5'b01111; w[53][184] = 5'b01111; w[53][185] = 5'b01111; w[53][186] = 5'b01111; w[53][187] = 5'b01111; w[53][188] = 5'b01111; w[53][189] = 5'b01111; w[53][190] = 5'b01111; w[53][191] = 5'b01111; w[53][192] = 5'b01111; w[53][193] = 5'b01111; w[53][194] = 5'b01111; w[53][195] = 5'b01111; w[53][196] = 5'b01111; w[53][197] = 5'b01111; w[53][198] = 5'b01111; w[53][199] = 5'b01111; w[53][200] = 5'b01111; w[53][201] = 5'b01111; w[53][202] = 5'b01111; w[53][203] = 5'b01111; w[53][204] = 5'b01111; w[53][205] = 5'b01111; w[53][206] = 5'b01111; w[53][207] = 5'b01111; w[53][208] = 5'b01111; w[53][209] = 5'b01111; 
w[54][0] = 5'b01111; w[54][1] = 5'b01111; w[54][2] = 5'b01111; w[54][3] = 5'b01111; w[54][4] = 5'b01111; w[54][5] = 5'b01111; w[54][6] = 5'b01111; w[54][7] = 5'b01111; w[54][8] = 5'b01111; w[54][9] = 5'b01111; w[54][10] = 5'b01111; w[54][11] = 5'b01111; w[54][12] = 5'b01111; w[54][13] = 5'b01111; w[54][14] = 5'b01111; w[54][15] = 5'b01111; w[54][16] = 5'b01111; w[54][17] = 5'b01111; w[54][18] = 5'b01111; w[54][19] = 5'b01111; w[54][20] = 5'b01111; w[54][21] = 5'b01111; w[54][22] = 5'b01111; w[54][23] = 5'b01111; w[54][24] = 5'b01111; w[54][25] = 5'b01111; w[54][26] = 5'b01111; w[54][27] = 5'b01111; w[54][28] = 5'b01111; w[54][29] = 5'b01111; w[54][30] = 5'b01111; w[54][31] = 5'b00000; w[54][32] = 5'b10000; w[54][33] = 5'b10000; w[54][34] = 5'b10000; w[54][35] = 5'b10000; w[54][36] = 5'b10000; w[54][37] = 5'b10000; w[54][38] = 5'b00000; w[54][39] = 5'b01111; w[54][40] = 5'b01111; w[54][41] = 5'b01111; w[54][42] = 5'b01111; w[54][43] = 5'b01111; w[54][44] = 5'b01111; w[54][45] = 5'b10000; w[54][46] = 5'b10000; w[54][47] = 5'b10000; w[54][48] = 5'b10000; w[54][49] = 5'b10000; w[54][50] = 5'b10000; w[54][51] = 5'b10000; w[54][52] = 5'b10000; w[54][53] = 5'b01111; w[54][54] = 5'b00000; w[54][55] = 5'b01111; w[54][56] = 5'b01111; w[54][57] = 5'b01111; w[54][58] = 5'b01111; w[54][59] = 5'b00000; w[54][60] = 5'b00000; w[54][61] = 5'b01111; w[54][62] = 5'b10000; w[54][63] = 5'b00000; w[54][64] = 5'b01111; w[54][65] = 5'b00000; w[54][66] = 5'b00000; w[54][67] = 5'b01111; w[54][68] = 5'b01111; w[54][69] = 5'b01111; w[54][70] = 5'b01111; w[54][71] = 5'b01111; w[54][72] = 5'b01111; w[54][73] = 5'b00000; w[54][74] = 5'b01111; w[54][75] = 5'b01111; w[54][76] = 5'b10000; w[54][77] = 5'b00000; w[54][78] = 5'b01111; w[54][79] = 5'b01111; w[54][80] = 5'b00000; w[54][81] = 5'b01111; w[54][82] = 5'b01111; w[54][83] = 5'b01111; w[54][84] = 5'b01111; w[54][85] = 5'b01111; w[54][86] = 5'b01111; w[54][87] = 5'b00000; w[54][88] = 5'b01111; w[54][89] = 5'b01111; w[54][90] = 5'b10000; w[54][91] = 5'b10000; w[54][92] = 5'b01111; w[54][93] = 5'b01111; w[54][94] = 5'b01111; w[54][95] = 5'b01111; w[54][96] = 5'b01111; w[54][97] = 5'b01111; w[54][98] = 5'b01111; w[54][99] = 5'b01111; w[54][100] = 5'b01111; w[54][101] = 5'b00000; w[54][102] = 5'b01111; w[54][103] = 5'b01111; w[54][104] = 5'b10000; w[54][105] = 5'b10000; w[54][106] = 5'b01111; w[54][107] = 5'b00000; w[54][108] = 5'b00000; w[54][109] = 5'b01111; w[54][110] = 5'b01111; w[54][111] = 5'b01111; w[54][112] = 5'b01111; w[54][113] = 5'b01111; w[54][114] = 5'b01111; w[54][115] = 5'b00000; w[54][116] = 5'b01111; w[54][117] = 5'b01111; w[54][118] = 5'b10000; w[54][119] = 5'b10000; w[54][120] = 5'b00000; w[54][121] = 5'b00000; w[54][122] = 5'b00000; w[54][123] = 5'b01111; w[54][124] = 5'b01111; w[54][125] = 5'b01111; w[54][126] = 5'b01111; w[54][127] = 5'b01111; w[54][128] = 5'b01111; w[54][129] = 5'b00000; w[54][130] = 5'b01111; w[54][131] = 5'b01111; w[54][132] = 5'b00000; w[54][133] = 5'b10000; w[54][134] = 5'b01111; w[54][135] = 5'b01111; w[54][136] = 5'b00000; w[54][137] = 5'b01111; w[54][138] = 5'b01111; w[54][139] = 5'b01111; w[54][140] = 5'b01111; w[54][141] = 5'b01111; w[54][142] = 5'b01111; w[54][143] = 5'b00000; w[54][144] = 5'b00000; w[54][145] = 5'b01111; w[54][146] = 5'b00000; w[54][147] = 5'b10000; w[54][148] = 5'b01111; w[54][149] = 5'b00000; w[54][150] = 5'b00000; w[54][151] = 5'b01111; w[54][152] = 5'b01111; w[54][153] = 5'b01111; w[54][154] = 5'b01111; w[54][155] = 5'b01111; w[54][156] = 5'b01111; w[54][157] = 5'b00000; w[54][158] = 5'b00000; w[54][159] = 5'b00000; w[54][160] = 5'b10000; w[54][161] = 5'b10000; w[54][162] = 5'b10000; w[54][163] = 5'b00000; w[54][164] = 5'b00000; w[54][165] = 5'b01111; w[54][166] = 5'b01111; w[54][167] = 5'b01111; w[54][168] = 5'b01111; w[54][169] = 5'b01111; w[54][170] = 5'b01111; w[54][171] = 5'b01111; w[54][172] = 5'b00000; w[54][173] = 5'b00000; w[54][174] = 5'b10000; w[54][175] = 5'b10000; w[54][176] = 5'b10000; w[54][177] = 5'b00000; w[54][178] = 5'b01111; w[54][179] = 5'b01111; w[54][180] = 5'b01111; w[54][181] = 5'b01111; w[54][182] = 5'b01111; w[54][183] = 5'b01111; w[54][184] = 5'b01111; w[54][185] = 5'b01111; w[54][186] = 5'b01111; w[54][187] = 5'b01111; w[54][188] = 5'b01111; w[54][189] = 5'b01111; w[54][190] = 5'b01111; w[54][191] = 5'b01111; w[54][192] = 5'b01111; w[54][193] = 5'b01111; w[54][194] = 5'b01111; w[54][195] = 5'b01111; w[54][196] = 5'b01111; w[54][197] = 5'b01111; w[54][198] = 5'b01111; w[54][199] = 5'b01111; w[54][200] = 5'b01111; w[54][201] = 5'b01111; w[54][202] = 5'b01111; w[54][203] = 5'b01111; w[54][204] = 5'b01111; w[54][205] = 5'b01111; w[54][206] = 5'b01111; w[54][207] = 5'b01111; w[54][208] = 5'b01111; w[54][209] = 5'b01111; 
w[55][0] = 5'b01111; w[55][1] = 5'b01111; w[55][2] = 5'b01111; w[55][3] = 5'b01111; w[55][4] = 5'b01111; w[55][5] = 5'b01111; w[55][6] = 5'b01111; w[55][7] = 5'b01111; w[55][8] = 5'b01111; w[55][9] = 5'b01111; w[55][10] = 5'b01111; w[55][11] = 5'b01111; w[55][12] = 5'b01111; w[55][13] = 5'b01111; w[55][14] = 5'b01111; w[55][15] = 5'b01111; w[55][16] = 5'b01111; w[55][17] = 5'b01111; w[55][18] = 5'b01111; w[55][19] = 5'b01111; w[55][20] = 5'b01111; w[55][21] = 5'b01111; w[55][22] = 5'b01111; w[55][23] = 5'b01111; w[55][24] = 5'b01111; w[55][25] = 5'b01111; w[55][26] = 5'b01111; w[55][27] = 5'b01111; w[55][28] = 5'b01111; w[55][29] = 5'b01111; w[55][30] = 5'b01111; w[55][31] = 5'b00000; w[55][32] = 5'b10000; w[55][33] = 5'b10000; w[55][34] = 5'b10000; w[55][35] = 5'b10000; w[55][36] = 5'b10000; w[55][37] = 5'b10000; w[55][38] = 5'b00000; w[55][39] = 5'b01111; w[55][40] = 5'b01111; w[55][41] = 5'b01111; w[55][42] = 5'b01111; w[55][43] = 5'b01111; w[55][44] = 5'b01111; w[55][45] = 5'b10000; w[55][46] = 5'b10000; w[55][47] = 5'b10000; w[55][48] = 5'b10000; w[55][49] = 5'b10000; w[55][50] = 5'b10000; w[55][51] = 5'b10000; w[55][52] = 5'b10000; w[55][53] = 5'b01111; w[55][54] = 5'b01111; w[55][55] = 5'b00000; w[55][56] = 5'b01111; w[55][57] = 5'b01111; w[55][58] = 5'b01111; w[55][59] = 5'b00000; w[55][60] = 5'b00000; w[55][61] = 5'b01111; w[55][62] = 5'b10000; w[55][63] = 5'b00000; w[55][64] = 5'b01111; w[55][65] = 5'b00000; w[55][66] = 5'b00000; w[55][67] = 5'b01111; w[55][68] = 5'b01111; w[55][69] = 5'b01111; w[55][70] = 5'b01111; w[55][71] = 5'b01111; w[55][72] = 5'b01111; w[55][73] = 5'b00000; w[55][74] = 5'b01111; w[55][75] = 5'b01111; w[55][76] = 5'b10000; w[55][77] = 5'b00000; w[55][78] = 5'b01111; w[55][79] = 5'b01111; w[55][80] = 5'b00000; w[55][81] = 5'b01111; w[55][82] = 5'b01111; w[55][83] = 5'b01111; w[55][84] = 5'b01111; w[55][85] = 5'b01111; w[55][86] = 5'b01111; w[55][87] = 5'b00000; w[55][88] = 5'b01111; w[55][89] = 5'b01111; w[55][90] = 5'b10000; w[55][91] = 5'b10000; w[55][92] = 5'b01111; w[55][93] = 5'b01111; w[55][94] = 5'b01111; w[55][95] = 5'b01111; w[55][96] = 5'b01111; w[55][97] = 5'b01111; w[55][98] = 5'b01111; w[55][99] = 5'b01111; w[55][100] = 5'b01111; w[55][101] = 5'b00000; w[55][102] = 5'b01111; w[55][103] = 5'b01111; w[55][104] = 5'b10000; w[55][105] = 5'b10000; w[55][106] = 5'b01111; w[55][107] = 5'b00000; w[55][108] = 5'b00000; w[55][109] = 5'b01111; w[55][110] = 5'b01111; w[55][111] = 5'b01111; w[55][112] = 5'b01111; w[55][113] = 5'b01111; w[55][114] = 5'b01111; w[55][115] = 5'b00000; w[55][116] = 5'b01111; w[55][117] = 5'b01111; w[55][118] = 5'b10000; w[55][119] = 5'b10000; w[55][120] = 5'b00000; w[55][121] = 5'b00000; w[55][122] = 5'b00000; w[55][123] = 5'b01111; w[55][124] = 5'b01111; w[55][125] = 5'b01111; w[55][126] = 5'b01111; w[55][127] = 5'b01111; w[55][128] = 5'b01111; w[55][129] = 5'b00000; w[55][130] = 5'b01111; w[55][131] = 5'b01111; w[55][132] = 5'b00000; w[55][133] = 5'b10000; w[55][134] = 5'b01111; w[55][135] = 5'b01111; w[55][136] = 5'b00000; w[55][137] = 5'b01111; w[55][138] = 5'b01111; w[55][139] = 5'b01111; w[55][140] = 5'b01111; w[55][141] = 5'b01111; w[55][142] = 5'b01111; w[55][143] = 5'b00000; w[55][144] = 5'b00000; w[55][145] = 5'b01111; w[55][146] = 5'b00000; w[55][147] = 5'b10000; w[55][148] = 5'b01111; w[55][149] = 5'b00000; w[55][150] = 5'b00000; w[55][151] = 5'b01111; w[55][152] = 5'b01111; w[55][153] = 5'b01111; w[55][154] = 5'b01111; w[55][155] = 5'b01111; w[55][156] = 5'b01111; w[55][157] = 5'b00000; w[55][158] = 5'b00000; w[55][159] = 5'b00000; w[55][160] = 5'b10000; w[55][161] = 5'b10000; w[55][162] = 5'b10000; w[55][163] = 5'b00000; w[55][164] = 5'b00000; w[55][165] = 5'b01111; w[55][166] = 5'b01111; w[55][167] = 5'b01111; w[55][168] = 5'b01111; w[55][169] = 5'b01111; w[55][170] = 5'b01111; w[55][171] = 5'b01111; w[55][172] = 5'b00000; w[55][173] = 5'b00000; w[55][174] = 5'b10000; w[55][175] = 5'b10000; w[55][176] = 5'b10000; w[55][177] = 5'b00000; w[55][178] = 5'b01111; w[55][179] = 5'b01111; w[55][180] = 5'b01111; w[55][181] = 5'b01111; w[55][182] = 5'b01111; w[55][183] = 5'b01111; w[55][184] = 5'b01111; w[55][185] = 5'b01111; w[55][186] = 5'b01111; w[55][187] = 5'b01111; w[55][188] = 5'b01111; w[55][189] = 5'b01111; w[55][190] = 5'b01111; w[55][191] = 5'b01111; w[55][192] = 5'b01111; w[55][193] = 5'b01111; w[55][194] = 5'b01111; w[55][195] = 5'b01111; w[55][196] = 5'b01111; w[55][197] = 5'b01111; w[55][198] = 5'b01111; w[55][199] = 5'b01111; w[55][200] = 5'b01111; w[55][201] = 5'b01111; w[55][202] = 5'b01111; w[55][203] = 5'b01111; w[55][204] = 5'b01111; w[55][205] = 5'b01111; w[55][206] = 5'b01111; w[55][207] = 5'b01111; w[55][208] = 5'b01111; w[55][209] = 5'b01111; 
w[56][0] = 5'b01111; w[56][1] = 5'b01111; w[56][2] = 5'b01111; w[56][3] = 5'b01111; w[56][4] = 5'b01111; w[56][5] = 5'b01111; w[56][6] = 5'b01111; w[56][7] = 5'b01111; w[56][8] = 5'b01111; w[56][9] = 5'b01111; w[56][10] = 5'b01111; w[56][11] = 5'b01111; w[56][12] = 5'b01111; w[56][13] = 5'b01111; w[56][14] = 5'b01111; w[56][15] = 5'b01111; w[56][16] = 5'b01111; w[56][17] = 5'b01111; w[56][18] = 5'b01111; w[56][19] = 5'b01111; w[56][20] = 5'b01111; w[56][21] = 5'b01111; w[56][22] = 5'b01111; w[56][23] = 5'b01111; w[56][24] = 5'b01111; w[56][25] = 5'b01111; w[56][26] = 5'b01111; w[56][27] = 5'b01111; w[56][28] = 5'b01111; w[56][29] = 5'b01111; w[56][30] = 5'b01111; w[56][31] = 5'b00000; w[56][32] = 5'b10000; w[56][33] = 5'b10000; w[56][34] = 5'b10000; w[56][35] = 5'b10000; w[56][36] = 5'b10000; w[56][37] = 5'b10000; w[56][38] = 5'b00000; w[56][39] = 5'b01111; w[56][40] = 5'b01111; w[56][41] = 5'b01111; w[56][42] = 5'b01111; w[56][43] = 5'b01111; w[56][44] = 5'b01111; w[56][45] = 5'b10000; w[56][46] = 5'b10000; w[56][47] = 5'b10000; w[56][48] = 5'b10000; w[56][49] = 5'b10000; w[56][50] = 5'b10000; w[56][51] = 5'b10000; w[56][52] = 5'b10000; w[56][53] = 5'b01111; w[56][54] = 5'b01111; w[56][55] = 5'b01111; w[56][56] = 5'b00000; w[56][57] = 5'b01111; w[56][58] = 5'b01111; w[56][59] = 5'b00000; w[56][60] = 5'b00000; w[56][61] = 5'b01111; w[56][62] = 5'b10000; w[56][63] = 5'b00000; w[56][64] = 5'b01111; w[56][65] = 5'b00000; w[56][66] = 5'b00000; w[56][67] = 5'b01111; w[56][68] = 5'b01111; w[56][69] = 5'b01111; w[56][70] = 5'b01111; w[56][71] = 5'b01111; w[56][72] = 5'b01111; w[56][73] = 5'b00000; w[56][74] = 5'b01111; w[56][75] = 5'b01111; w[56][76] = 5'b10000; w[56][77] = 5'b00000; w[56][78] = 5'b01111; w[56][79] = 5'b01111; w[56][80] = 5'b00000; w[56][81] = 5'b01111; w[56][82] = 5'b01111; w[56][83] = 5'b01111; w[56][84] = 5'b01111; w[56][85] = 5'b01111; w[56][86] = 5'b01111; w[56][87] = 5'b00000; w[56][88] = 5'b01111; w[56][89] = 5'b01111; w[56][90] = 5'b10000; w[56][91] = 5'b10000; w[56][92] = 5'b01111; w[56][93] = 5'b01111; w[56][94] = 5'b01111; w[56][95] = 5'b01111; w[56][96] = 5'b01111; w[56][97] = 5'b01111; w[56][98] = 5'b01111; w[56][99] = 5'b01111; w[56][100] = 5'b01111; w[56][101] = 5'b00000; w[56][102] = 5'b01111; w[56][103] = 5'b01111; w[56][104] = 5'b10000; w[56][105] = 5'b10000; w[56][106] = 5'b01111; w[56][107] = 5'b00000; w[56][108] = 5'b00000; w[56][109] = 5'b01111; w[56][110] = 5'b01111; w[56][111] = 5'b01111; w[56][112] = 5'b01111; w[56][113] = 5'b01111; w[56][114] = 5'b01111; w[56][115] = 5'b00000; w[56][116] = 5'b01111; w[56][117] = 5'b01111; w[56][118] = 5'b10000; w[56][119] = 5'b10000; w[56][120] = 5'b00000; w[56][121] = 5'b00000; w[56][122] = 5'b00000; w[56][123] = 5'b01111; w[56][124] = 5'b01111; w[56][125] = 5'b01111; w[56][126] = 5'b01111; w[56][127] = 5'b01111; w[56][128] = 5'b01111; w[56][129] = 5'b00000; w[56][130] = 5'b01111; w[56][131] = 5'b01111; w[56][132] = 5'b00000; w[56][133] = 5'b10000; w[56][134] = 5'b01111; w[56][135] = 5'b01111; w[56][136] = 5'b00000; w[56][137] = 5'b01111; w[56][138] = 5'b01111; w[56][139] = 5'b01111; w[56][140] = 5'b01111; w[56][141] = 5'b01111; w[56][142] = 5'b01111; w[56][143] = 5'b00000; w[56][144] = 5'b00000; w[56][145] = 5'b01111; w[56][146] = 5'b00000; w[56][147] = 5'b10000; w[56][148] = 5'b01111; w[56][149] = 5'b00000; w[56][150] = 5'b00000; w[56][151] = 5'b01111; w[56][152] = 5'b01111; w[56][153] = 5'b01111; w[56][154] = 5'b01111; w[56][155] = 5'b01111; w[56][156] = 5'b01111; w[56][157] = 5'b00000; w[56][158] = 5'b00000; w[56][159] = 5'b00000; w[56][160] = 5'b10000; w[56][161] = 5'b10000; w[56][162] = 5'b10000; w[56][163] = 5'b00000; w[56][164] = 5'b00000; w[56][165] = 5'b01111; w[56][166] = 5'b01111; w[56][167] = 5'b01111; w[56][168] = 5'b01111; w[56][169] = 5'b01111; w[56][170] = 5'b01111; w[56][171] = 5'b01111; w[56][172] = 5'b00000; w[56][173] = 5'b00000; w[56][174] = 5'b10000; w[56][175] = 5'b10000; w[56][176] = 5'b10000; w[56][177] = 5'b00000; w[56][178] = 5'b01111; w[56][179] = 5'b01111; w[56][180] = 5'b01111; w[56][181] = 5'b01111; w[56][182] = 5'b01111; w[56][183] = 5'b01111; w[56][184] = 5'b01111; w[56][185] = 5'b01111; w[56][186] = 5'b01111; w[56][187] = 5'b01111; w[56][188] = 5'b01111; w[56][189] = 5'b01111; w[56][190] = 5'b01111; w[56][191] = 5'b01111; w[56][192] = 5'b01111; w[56][193] = 5'b01111; w[56][194] = 5'b01111; w[56][195] = 5'b01111; w[56][196] = 5'b01111; w[56][197] = 5'b01111; w[56][198] = 5'b01111; w[56][199] = 5'b01111; w[56][200] = 5'b01111; w[56][201] = 5'b01111; w[56][202] = 5'b01111; w[56][203] = 5'b01111; w[56][204] = 5'b01111; w[56][205] = 5'b01111; w[56][206] = 5'b01111; w[56][207] = 5'b01111; w[56][208] = 5'b01111; w[56][209] = 5'b01111; 
w[57][0] = 5'b01111; w[57][1] = 5'b01111; w[57][2] = 5'b01111; w[57][3] = 5'b01111; w[57][4] = 5'b01111; w[57][5] = 5'b01111; w[57][6] = 5'b01111; w[57][7] = 5'b01111; w[57][8] = 5'b01111; w[57][9] = 5'b01111; w[57][10] = 5'b01111; w[57][11] = 5'b01111; w[57][12] = 5'b01111; w[57][13] = 5'b01111; w[57][14] = 5'b01111; w[57][15] = 5'b01111; w[57][16] = 5'b01111; w[57][17] = 5'b01111; w[57][18] = 5'b01111; w[57][19] = 5'b01111; w[57][20] = 5'b01111; w[57][21] = 5'b01111; w[57][22] = 5'b01111; w[57][23] = 5'b01111; w[57][24] = 5'b01111; w[57][25] = 5'b01111; w[57][26] = 5'b01111; w[57][27] = 5'b01111; w[57][28] = 5'b01111; w[57][29] = 5'b01111; w[57][30] = 5'b01111; w[57][31] = 5'b00000; w[57][32] = 5'b10000; w[57][33] = 5'b10000; w[57][34] = 5'b10000; w[57][35] = 5'b10000; w[57][36] = 5'b10000; w[57][37] = 5'b10000; w[57][38] = 5'b00000; w[57][39] = 5'b01111; w[57][40] = 5'b01111; w[57][41] = 5'b01111; w[57][42] = 5'b01111; w[57][43] = 5'b01111; w[57][44] = 5'b01111; w[57][45] = 5'b10000; w[57][46] = 5'b10000; w[57][47] = 5'b10000; w[57][48] = 5'b10000; w[57][49] = 5'b10000; w[57][50] = 5'b10000; w[57][51] = 5'b10000; w[57][52] = 5'b10000; w[57][53] = 5'b01111; w[57][54] = 5'b01111; w[57][55] = 5'b01111; w[57][56] = 5'b01111; w[57][57] = 5'b00000; w[57][58] = 5'b01111; w[57][59] = 5'b00000; w[57][60] = 5'b00000; w[57][61] = 5'b01111; w[57][62] = 5'b10000; w[57][63] = 5'b00000; w[57][64] = 5'b01111; w[57][65] = 5'b00000; w[57][66] = 5'b00000; w[57][67] = 5'b01111; w[57][68] = 5'b01111; w[57][69] = 5'b01111; w[57][70] = 5'b01111; w[57][71] = 5'b01111; w[57][72] = 5'b01111; w[57][73] = 5'b00000; w[57][74] = 5'b01111; w[57][75] = 5'b01111; w[57][76] = 5'b10000; w[57][77] = 5'b00000; w[57][78] = 5'b01111; w[57][79] = 5'b01111; w[57][80] = 5'b00000; w[57][81] = 5'b01111; w[57][82] = 5'b01111; w[57][83] = 5'b01111; w[57][84] = 5'b01111; w[57][85] = 5'b01111; w[57][86] = 5'b01111; w[57][87] = 5'b00000; w[57][88] = 5'b01111; w[57][89] = 5'b01111; w[57][90] = 5'b10000; w[57][91] = 5'b10000; w[57][92] = 5'b01111; w[57][93] = 5'b01111; w[57][94] = 5'b01111; w[57][95] = 5'b01111; w[57][96] = 5'b01111; w[57][97] = 5'b01111; w[57][98] = 5'b01111; w[57][99] = 5'b01111; w[57][100] = 5'b01111; w[57][101] = 5'b00000; w[57][102] = 5'b01111; w[57][103] = 5'b01111; w[57][104] = 5'b10000; w[57][105] = 5'b10000; w[57][106] = 5'b01111; w[57][107] = 5'b00000; w[57][108] = 5'b00000; w[57][109] = 5'b01111; w[57][110] = 5'b01111; w[57][111] = 5'b01111; w[57][112] = 5'b01111; w[57][113] = 5'b01111; w[57][114] = 5'b01111; w[57][115] = 5'b00000; w[57][116] = 5'b01111; w[57][117] = 5'b01111; w[57][118] = 5'b10000; w[57][119] = 5'b10000; w[57][120] = 5'b00000; w[57][121] = 5'b00000; w[57][122] = 5'b00000; w[57][123] = 5'b01111; w[57][124] = 5'b01111; w[57][125] = 5'b01111; w[57][126] = 5'b01111; w[57][127] = 5'b01111; w[57][128] = 5'b01111; w[57][129] = 5'b00000; w[57][130] = 5'b01111; w[57][131] = 5'b01111; w[57][132] = 5'b00000; w[57][133] = 5'b10000; w[57][134] = 5'b01111; w[57][135] = 5'b01111; w[57][136] = 5'b00000; w[57][137] = 5'b01111; w[57][138] = 5'b01111; w[57][139] = 5'b01111; w[57][140] = 5'b01111; w[57][141] = 5'b01111; w[57][142] = 5'b01111; w[57][143] = 5'b00000; w[57][144] = 5'b00000; w[57][145] = 5'b01111; w[57][146] = 5'b00000; w[57][147] = 5'b10000; w[57][148] = 5'b01111; w[57][149] = 5'b00000; w[57][150] = 5'b00000; w[57][151] = 5'b01111; w[57][152] = 5'b01111; w[57][153] = 5'b01111; w[57][154] = 5'b01111; w[57][155] = 5'b01111; w[57][156] = 5'b01111; w[57][157] = 5'b00000; w[57][158] = 5'b00000; w[57][159] = 5'b00000; w[57][160] = 5'b10000; w[57][161] = 5'b10000; w[57][162] = 5'b10000; w[57][163] = 5'b00000; w[57][164] = 5'b00000; w[57][165] = 5'b01111; w[57][166] = 5'b01111; w[57][167] = 5'b01111; w[57][168] = 5'b01111; w[57][169] = 5'b01111; w[57][170] = 5'b01111; w[57][171] = 5'b01111; w[57][172] = 5'b00000; w[57][173] = 5'b00000; w[57][174] = 5'b10000; w[57][175] = 5'b10000; w[57][176] = 5'b10000; w[57][177] = 5'b00000; w[57][178] = 5'b01111; w[57][179] = 5'b01111; w[57][180] = 5'b01111; w[57][181] = 5'b01111; w[57][182] = 5'b01111; w[57][183] = 5'b01111; w[57][184] = 5'b01111; w[57][185] = 5'b01111; w[57][186] = 5'b01111; w[57][187] = 5'b01111; w[57][188] = 5'b01111; w[57][189] = 5'b01111; w[57][190] = 5'b01111; w[57][191] = 5'b01111; w[57][192] = 5'b01111; w[57][193] = 5'b01111; w[57][194] = 5'b01111; w[57][195] = 5'b01111; w[57][196] = 5'b01111; w[57][197] = 5'b01111; w[57][198] = 5'b01111; w[57][199] = 5'b01111; w[57][200] = 5'b01111; w[57][201] = 5'b01111; w[57][202] = 5'b01111; w[57][203] = 5'b01111; w[57][204] = 5'b01111; w[57][205] = 5'b01111; w[57][206] = 5'b01111; w[57][207] = 5'b01111; w[57][208] = 5'b01111; w[57][209] = 5'b01111; 
w[58][0] = 5'b01111; w[58][1] = 5'b01111; w[58][2] = 5'b01111; w[58][3] = 5'b01111; w[58][4] = 5'b01111; w[58][5] = 5'b01111; w[58][6] = 5'b01111; w[58][7] = 5'b01111; w[58][8] = 5'b01111; w[58][9] = 5'b01111; w[58][10] = 5'b01111; w[58][11] = 5'b01111; w[58][12] = 5'b01111; w[58][13] = 5'b01111; w[58][14] = 5'b01111; w[58][15] = 5'b01111; w[58][16] = 5'b01111; w[58][17] = 5'b01111; w[58][18] = 5'b01111; w[58][19] = 5'b01111; w[58][20] = 5'b01111; w[58][21] = 5'b01111; w[58][22] = 5'b01111; w[58][23] = 5'b01111; w[58][24] = 5'b01111; w[58][25] = 5'b01111; w[58][26] = 5'b01111; w[58][27] = 5'b01111; w[58][28] = 5'b01111; w[58][29] = 5'b01111; w[58][30] = 5'b00000; w[58][31] = 5'b10000; w[58][32] = 5'b00000; w[58][33] = 5'b10000; w[58][34] = 5'b00000; w[58][35] = 5'b00000; w[58][36] = 5'b00000; w[58][37] = 5'b00000; w[58][38] = 5'b10000; w[58][39] = 5'b00000; w[58][40] = 5'b01111; w[58][41] = 5'b01111; w[58][42] = 5'b01111; w[58][43] = 5'b01111; w[58][44] = 5'b00000; w[58][45] = 5'b00000; w[58][46] = 5'b00000; w[58][47] = 5'b10000; w[58][48] = 5'b00000; w[58][49] = 5'b00000; w[58][50] = 5'b00000; w[58][51] = 5'b00000; w[58][52] = 5'b00000; w[58][53] = 5'b00000; w[58][54] = 5'b01111; w[58][55] = 5'b01111; w[58][56] = 5'b01111; w[58][57] = 5'b01111; w[58][58] = 5'b00000; w[58][59] = 5'b01111; w[58][60] = 5'b01111; w[58][61] = 5'b00000; w[58][62] = 5'b10000; w[58][63] = 5'b10000; w[58][64] = 5'b01111; w[58][65] = 5'b01111; w[58][66] = 5'b01111; w[58][67] = 5'b01111; w[58][68] = 5'b01111; w[58][69] = 5'b01111; w[58][70] = 5'b01111; w[58][71] = 5'b01111; w[58][72] = 5'b01111; w[58][73] = 5'b01111; w[58][74] = 5'b00000; w[58][75] = 5'b00000; w[58][76] = 5'b10000; w[58][77] = 5'b10000; w[58][78] = 5'b01111; w[58][79] = 5'b00000; w[58][80] = 5'b01111; w[58][81] = 5'b01111; w[58][82] = 5'b01111; w[58][83] = 5'b01111; w[58][84] = 5'b01111; w[58][85] = 5'b01111; w[58][86] = 5'b01111; w[58][87] = 5'b01111; w[58][88] = 5'b00000; w[58][89] = 5'b00000; w[58][90] = 5'b10000; w[58][91] = 5'b10000; w[58][92] = 5'b01111; w[58][93] = 5'b00000; w[58][94] = 5'b00000; w[58][95] = 5'b01111; w[58][96] = 5'b01111; w[58][97] = 5'b01111; w[58][98] = 5'b01111; w[58][99] = 5'b01111; w[58][100] = 5'b01111; w[58][101] = 5'b01111; w[58][102] = 5'b00000; w[58][103] = 5'b01111; w[58][104] = 5'b10000; w[58][105] = 5'b10000; w[58][106] = 5'b01111; w[58][107] = 5'b01111; w[58][108] = 5'b01111; w[58][109] = 5'b01111; w[58][110] = 5'b01111; w[58][111] = 5'b01111; w[58][112] = 5'b01111; w[58][113] = 5'b01111; w[58][114] = 5'b01111; w[58][115] = 5'b01111; w[58][116] = 5'b00000; w[58][117] = 5'b01111; w[58][118] = 5'b10000; w[58][119] = 5'b10000; w[58][120] = 5'b01111; w[58][121] = 5'b01111; w[58][122] = 5'b01111; w[58][123] = 5'b01111; w[58][124] = 5'b01111; w[58][125] = 5'b01111; w[58][126] = 5'b01111; w[58][127] = 5'b01111; w[58][128] = 5'b01111; w[58][129] = 5'b01111; w[58][130] = 5'b00000; w[58][131] = 5'b01111; w[58][132] = 5'b10000; w[58][133] = 5'b10000; w[58][134] = 5'b00000; w[58][135] = 5'b00000; w[58][136] = 5'b01111; w[58][137] = 5'b01111; w[58][138] = 5'b01111; w[58][139] = 5'b01111; w[58][140] = 5'b01111; w[58][141] = 5'b01111; w[58][142] = 5'b01111; w[58][143] = 5'b01111; w[58][144] = 5'b01111; w[58][145] = 5'b01111; w[58][146] = 5'b10000; w[58][147] = 5'b10000; w[58][148] = 5'b00000; w[58][149] = 5'b01111; w[58][150] = 5'b01111; w[58][151] = 5'b01111; w[58][152] = 5'b01111; w[58][153] = 5'b01111; w[58][154] = 5'b01111; w[58][155] = 5'b01111; w[58][156] = 5'b01111; w[58][157] = 5'b01111; w[58][158] = 5'b01111; w[58][159] = 5'b01111; w[58][160] = 5'b00000; w[58][161] = 5'b00000; w[58][162] = 5'b00000; w[58][163] = 5'b01111; w[58][164] = 5'b01111; w[58][165] = 5'b01111; w[58][166] = 5'b01111; w[58][167] = 5'b01111; w[58][168] = 5'b01111; w[58][169] = 5'b01111; w[58][170] = 5'b01111; w[58][171] = 5'b00000; w[58][172] = 5'b01111; w[58][173] = 5'b01111; w[58][174] = 5'b00000; w[58][175] = 5'b00000; w[58][176] = 5'b00000; w[58][177] = 5'b01111; w[58][178] = 5'b00000; w[58][179] = 5'b01111; w[58][180] = 5'b01111; w[58][181] = 5'b01111; w[58][182] = 5'b01111; w[58][183] = 5'b01111; w[58][184] = 5'b01111; w[58][185] = 5'b01111; w[58][186] = 5'b01111; w[58][187] = 5'b01111; w[58][188] = 5'b01111; w[58][189] = 5'b01111; w[58][190] = 5'b01111; w[58][191] = 5'b01111; w[58][192] = 5'b01111; w[58][193] = 5'b01111; w[58][194] = 5'b01111; w[58][195] = 5'b01111; w[58][196] = 5'b01111; w[58][197] = 5'b01111; w[58][198] = 5'b01111; w[58][199] = 5'b01111; w[58][200] = 5'b01111; w[58][201] = 5'b01111; w[58][202] = 5'b01111; w[58][203] = 5'b01111; w[58][204] = 5'b01111; w[58][205] = 5'b01111; w[58][206] = 5'b01111; w[58][207] = 5'b01111; w[58][208] = 5'b01111; w[58][209] = 5'b01111; 
w[59][0] = 5'b00000; w[59][1] = 5'b00000; w[59][2] = 5'b00000; w[59][3] = 5'b00000; w[59][4] = 5'b00000; w[59][5] = 5'b00000; w[59][6] = 5'b00000; w[59][7] = 5'b00000; w[59][8] = 5'b00000; w[59][9] = 5'b00000; w[59][10] = 5'b00000; w[59][11] = 5'b00000; w[59][12] = 5'b00000; w[59][13] = 5'b00000; w[59][14] = 5'b00000; w[59][15] = 5'b00000; w[59][16] = 5'b00000; w[59][17] = 5'b00000; w[59][18] = 5'b00000; w[59][19] = 5'b00000; w[59][20] = 5'b00000; w[59][21] = 5'b00000; w[59][22] = 5'b00000; w[59][23] = 5'b00000; w[59][24] = 5'b00000; w[59][25] = 5'b00000; w[59][26] = 5'b00000; w[59][27] = 5'b00000; w[59][28] = 5'b00000; w[59][29] = 5'b00000; w[59][30] = 5'b10000; w[59][31] = 5'b00000; w[59][32] = 5'b01111; w[59][33] = 5'b00000; w[59][34] = 5'b10000; w[59][35] = 5'b10000; w[59][36] = 5'b10000; w[59][37] = 5'b01111; w[59][38] = 5'b00000; w[59][39] = 5'b10000; w[59][40] = 5'b00000; w[59][41] = 5'b00000; w[59][42] = 5'b00000; w[59][43] = 5'b00000; w[59][44] = 5'b10000; w[59][45] = 5'b01111; w[59][46] = 5'b01111; w[59][47] = 5'b00000; w[59][48] = 5'b10000; w[59][49] = 5'b10000; w[59][50] = 5'b10000; w[59][51] = 5'b01111; w[59][52] = 5'b01111; w[59][53] = 5'b10000; w[59][54] = 5'b00000; w[59][55] = 5'b00000; w[59][56] = 5'b00000; w[59][57] = 5'b00000; w[59][58] = 5'b01111; w[59][59] = 5'b00000; w[59][60] = 5'b01111; w[59][61] = 5'b01111; w[59][62] = 5'b10000; w[59][63] = 5'b10000; w[59][64] = 5'b00000; w[59][65] = 5'b01111; w[59][66] = 5'b01111; w[59][67] = 5'b01111; w[59][68] = 5'b00000; w[59][69] = 5'b00000; w[59][70] = 5'b00000; w[59][71] = 5'b00000; w[59][72] = 5'b01111; w[59][73] = 5'b01111; w[59][74] = 5'b01111; w[59][75] = 5'b01111; w[59][76] = 5'b10000; w[59][77] = 5'b10000; w[59][78] = 5'b00000; w[59][79] = 5'b01111; w[59][80] = 5'b01111; w[59][81] = 5'b01111; w[59][82] = 5'b00000; w[59][83] = 5'b00000; w[59][84] = 5'b00000; w[59][85] = 5'b00000; w[59][86] = 5'b01111; w[59][87] = 5'b01111; w[59][88] = 5'b01111; w[59][89] = 5'b01111; w[59][90] = 5'b10000; w[59][91] = 5'b10000; w[59][92] = 5'b00000; w[59][93] = 5'b01111; w[59][94] = 5'b01111; w[59][95] = 5'b00000; w[59][96] = 5'b00000; w[59][97] = 5'b00000; w[59][98] = 5'b00000; w[59][99] = 5'b00000; w[59][100] = 5'b01111; w[59][101] = 5'b01111; w[59][102] = 5'b01111; w[59][103] = 5'b00000; w[59][104] = 5'b10000; w[59][105] = 5'b10000; w[59][106] = 5'b01111; w[59][107] = 5'b01111; w[59][108] = 5'b01111; w[59][109] = 5'b01111; w[59][110] = 5'b00000; w[59][111] = 5'b00000; w[59][112] = 5'b00000; w[59][113] = 5'b00000; w[59][114] = 5'b01111; w[59][115] = 5'b01111; w[59][116] = 5'b01111; w[59][117] = 5'b00000; w[59][118] = 5'b10000; w[59][119] = 5'b10000; w[59][120] = 5'b01111; w[59][121] = 5'b01111; w[59][122] = 5'b01111; w[59][123] = 5'b01111; w[59][124] = 5'b00000; w[59][125] = 5'b00000; w[59][126] = 5'b00000; w[59][127] = 5'b00000; w[59][128] = 5'b01111; w[59][129] = 5'b01111; w[59][130] = 5'b01111; w[59][131] = 5'b00000; w[59][132] = 5'b10000; w[59][133] = 5'b10000; w[59][134] = 5'b01111; w[59][135] = 5'b01111; w[59][136] = 5'b01111; w[59][137] = 5'b01111; w[59][138] = 5'b00000; w[59][139] = 5'b00000; w[59][140] = 5'b00000; w[59][141] = 5'b00000; w[59][142] = 5'b01111; w[59][143] = 5'b01111; w[59][144] = 5'b01111; w[59][145] = 5'b00000; w[59][146] = 5'b10000; w[59][147] = 5'b10000; w[59][148] = 5'b01111; w[59][149] = 5'b01111; w[59][150] = 5'b01111; w[59][151] = 5'b01111; w[59][152] = 5'b00000; w[59][153] = 5'b00000; w[59][154] = 5'b00000; w[59][155] = 5'b00000; w[59][156] = 5'b00000; w[59][157] = 5'b01111; w[59][158] = 5'b01111; w[59][159] = 5'b00000; w[59][160] = 5'b10000; w[59][161] = 5'b10000; w[59][162] = 5'b01111; w[59][163] = 5'b01111; w[59][164] = 5'b01111; w[59][165] = 5'b00000; w[59][166] = 5'b00000; w[59][167] = 5'b00000; w[59][168] = 5'b00000; w[59][169] = 5'b00000; w[59][170] = 5'b00000; w[59][171] = 5'b01111; w[59][172] = 5'b01111; w[59][173] = 5'b00000; w[59][174] = 5'b10000; w[59][175] = 5'b10000; w[59][176] = 5'b01111; w[59][177] = 5'b01111; w[59][178] = 5'b01111; w[59][179] = 5'b00000; w[59][180] = 5'b00000; w[59][181] = 5'b00000; w[59][182] = 5'b00000; w[59][183] = 5'b00000; w[59][184] = 5'b00000; w[59][185] = 5'b00000; w[59][186] = 5'b00000; w[59][187] = 5'b00000; w[59][188] = 5'b00000; w[59][189] = 5'b00000; w[59][190] = 5'b00000; w[59][191] = 5'b00000; w[59][192] = 5'b00000; w[59][193] = 5'b00000; w[59][194] = 5'b00000; w[59][195] = 5'b00000; w[59][196] = 5'b00000; w[59][197] = 5'b00000; w[59][198] = 5'b00000; w[59][199] = 5'b00000; w[59][200] = 5'b00000; w[59][201] = 5'b00000; w[59][202] = 5'b00000; w[59][203] = 5'b00000; w[59][204] = 5'b00000; w[59][205] = 5'b00000; w[59][206] = 5'b00000; w[59][207] = 5'b00000; w[59][208] = 5'b00000; w[59][209] = 5'b00000; 
w[60][0] = 5'b00000; w[60][1] = 5'b00000; w[60][2] = 5'b00000; w[60][3] = 5'b00000; w[60][4] = 5'b00000; w[60][5] = 5'b00000; w[60][6] = 5'b00000; w[60][7] = 5'b00000; w[60][8] = 5'b00000; w[60][9] = 5'b00000; w[60][10] = 5'b00000; w[60][11] = 5'b00000; w[60][12] = 5'b00000; w[60][13] = 5'b00000; w[60][14] = 5'b00000; w[60][15] = 5'b00000; w[60][16] = 5'b00000; w[60][17] = 5'b00000; w[60][18] = 5'b00000; w[60][19] = 5'b00000; w[60][20] = 5'b00000; w[60][21] = 5'b00000; w[60][22] = 5'b00000; w[60][23] = 5'b00000; w[60][24] = 5'b00000; w[60][25] = 5'b00000; w[60][26] = 5'b00000; w[60][27] = 5'b00000; w[60][28] = 5'b00000; w[60][29] = 5'b00000; w[60][30] = 5'b10000; w[60][31] = 5'b00000; w[60][32] = 5'b01111; w[60][33] = 5'b00000; w[60][34] = 5'b10000; w[60][35] = 5'b10000; w[60][36] = 5'b10000; w[60][37] = 5'b01111; w[60][38] = 5'b00000; w[60][39] = 5'b10000; w[60][40] = 5'b00000; w[60][41] = 5'b00000; w[60][42] = 5'b00000; w[60][43] = 5'b00000; w[60][44] = 5'b10000; w[60][45] = 5'b01111; w[60][46] = 5'b01111; w[60][47] = 5'b00000; w[60][48] = 5'b10000; w[60][49] = 5'b10000; w[60][50] = 5'b10000; w[60][51] = 5'b01111; w[60][52] = 5'b01111; w[60][53] = 5'b10000; w[60][54] = 5'b00000; w[60][55] = 5'b00000; w[60][56] = 5'b00000; w[60][57] = 5'b00000; w[60][58] = 5'b01111; w[60][59] = 5'b01111; w[60][60] = 5'b00000; w[60][61] = 5'b01111; w[60][62] = 5'b10000; w[60][63] = 5'b10000; w[60][64] = 5'b00000; w[60][65] = 5'b01111; w[60][66] = 5'b01111; w[60][67] = 5'b01111; w[60][68] = 5'b00000; w[60][69] = 5'b00000; w[60][70] = 5'b00000; w[60][71] = 5'b00000; w[60][72] = 5'b01111; w[60][73] = 5'b01111; w[60][74] = 5'b01111; w[60][75] = 5'b01111; w[60][76] = 5'b10000; w[60][77] = 5'b10000; w[60][78] = 5'b00000; w[60][79] = 5'b01111; w[60][80] = 5'b01111; w[60][81] = 5'b01111; w[60][82] = 5'b00000; w[60][83] = 5'b00000; w[60][84] = 5'b00000; w[60][85] = 5'b00000; w[60][86] = 5'b01111; w[60][87] = 5'b01111; w[60][88] = 5'b01111; w[60][89] = 5'b01111; w[60][90] = 5'b10000; w[60][91] = 5'b10000; w[60][92] = 5'b00000; w[60][93] = 5'b01111; w[60][94] = 5'b01111; w[60][95] = 5'b00000; w[60][96] = 5'b00000; w[60][97] = 5'b00000; w[60][98] = 5'b00000; w[60][99] = 5'b00000; w[60][100] = 5'b01111; w[60][101] = 5'b01111; w[60][102] = 5'b01111; w[60][103] = 5'b00000; w[60][104] = 5'b10000; w[60][105] = 5'b10000; w[60][106] = 5'b01111; w[60][107] = 5'b01111; w[60][108] = 5'b01111; w[60][109] = 5'b01111; w[60][110] = 5'b00000; w[60][111] = 5'b00000; w[60][112] = 5'b00000; w[60][113] = 5'b00000; w[60][114] = 5'b01111; w[60][115] = 5'b01111; w[60][116] = 5'b01111; w[60][117] = 5'b00000; w[60][118] = 5'b10000; w[60][119] = 5'b10000; w[60][120] = 5'b01111; w[60][121] = 5'b01111; w[60][122] = 5'b01111; w[60][123] = 5'b01111; w[60][124] = 5'b00000; w[60][125] = 5'b00000; w[60][126] = 5'b00000; w[60][127] = 5'b00000; w[60][128] = 5'b01111; w[60][129] = 5'b01111; w[60][130] = 5'b01111; w[60][131] = 5'b00000; w[60][132] = 5'b10000; w[60][133] = 5'b10000; w[60][134] = 5'b01111; w[60][135] = 5'b01111; w[60][136] = 5'b01111; w[60][137] = 5'b01111; w[60][138] = 5'b00000; w[60][139] = 5'b00000; w[60][140] = 5'b00000; w[60][141] = 5'b00000; w[60][142] = 5'b01111; w[60][143] = 5'b01111; w[60][144] = 5'b01111; w[60][145] = 5'b00000; w[60][146] = 5'b10000; w[60][147] = 5'b10000; w[60][148] = 5'b01111; w[60][149] = 5'b01111; w[60][150] = 5'b01111; w[60][151] = 5'b01111; w[60][152] = 5'b00000; w[60][153] = 5'b00000; w[60][154] = 5'b00000; w[60][155] = 5'b00000; w[60][156] = 5'b00000; w[60][157] = 5'b01111; w[60][158] = 5'b01111; w[60][159] = 5'b00000; w[60][160] = 5'b10000; w[60][161] = 5'b10000; w[60][162] = 5'b01111; w[60][163] = 5'b01111; w[60][164] = 5'b01111; w[60][165] = 5'b00000; w[60][166] = 5'b00000; w[60][167] = 5'b00000; w[60][168] = 5'b00000; w[60][169] = 5'b00000; w[60][170] = 5'b00000; w[60][171] = 5'b01111; w[60][172] = 5'b01111; w[60][173] = 5'b00000; w[60][174] = 5'b10000; w[60][175] = 5'b10000; w[60][176] = 5'b01111; w[60][177] = 5'b01111; w[60][178] = 5'b01111; w[60][179] = 5'b00000; w[60][180] = 5'b00000; w[60][181] = 5'b00000; w[60][182] = 5'b00000; w[60][183] = 5'b00000; w[60][184] = 5'b00000; w[60][185] = 5'b00000; w[60][186] = 5'b00000; w[60][187] = 5'b00000; w[60][188] = 5'b00000; w[60][189] = 5'b00000; w[60][190] = 5'b00000; w[60][191] = 5'b00000; w[60][192] = 5'b00000; w[60][193] = 5'b00000; w[60][194] = 5'b00000; w[60][195] = 5'b00000; w[60][196] = 5'b00000; w[60][197] = 5'b00000; w[60][198] = 5'b00000; w[60][199] = 5'b00000; w[60][200] = 5'b00000; w[60][201] = 5'b00000; w[60][202] = 5'b00000; w[60][203] = 5'b00000; w[60][204] = 5'b00000; w[60][205] = 5'b00000; w[60][206] = 5'b00000; w[60][207] = 5'b00000; w[60][208] = 5'b00000; w[60][209] = 5'b00000; 
w[61][0] = 5'b01111; w[61][1] = 5'b01111; w[61][2] = 5'b01111; w[61][3] = 5'b01111; w[61][4] = 5'b01111; w[61][5] = 5'b01111; w[61][6] = 5'b01111; w[61][7] = 5'b01111; w[61][8] = 5'b01111; w[61][9] = 5'b01111; w[61][10] = 5'b01111; w[61][11] = 5'b01111; w[61][12] = 5'b01111; w[61][13] = 5'b01111; w[61][14] = 5'b01111; w[61][15] = 5'b01111; w[61][16] = 5'b01111; w[61][17] = 5'b01111; w[61][18] = 5'b01111; w[61][19] = 5'b01111; w[61][20] = 5'b01111; w[61][21] = 5'b01111; w[61][22] = 5'b01111; w[61][23] = 5'b01111; w[61][24] = 5'b01111; w[61][25] = 5'b01111; w[61][26] = 5'b01111; w[61][27] = 5'b01111; w[61][28] = 5'b01111; w[61][29] = 5'b01111; w[61][30] = 5'b00000; w[61][31] = 5'b01111; w[61][32] = 5'b00000; w[61][33] = 5'b10000; w[61][34] = 5'b10000; w[61][35] = 5'b10000; w[61][36] = 5'b10000; w[61][37] = 5'b00000; w[61][38] = 5'b01111; w[61][39] = 5'b00000; w[61][40] = 5'b01111; w[61][41] = 5'b01111; w[61][42] = 5'b01111; w[61][43] = 5'b01111; w[61][44] = 5'b00000; w[61][45] = 5'b00000; w[61][46] = 5'b00000; w[61][47] = 5'b10000; w[61][48] = 5'b10000; w[61][49] = 5'b10000; w[61][50] = 5'b10000; w[61][51] = 5'b00000; w[61][52] = 5'b00000; w[61][53] = 5'b00000; w[61][54] = 5'b01111; w[61][55] = 5'b01111; w[61][56] = 5'b01111; w[61][57] = 5'b01111; w[61][58] = 5'b00000; w[61][59] = 5'b01111; w[61][60] = 5'b01111; w[61][61] = 5'b00000; w[61][62] = 5'b00000; w[61][63] = 5'b10000; w[61][64] = 5'b01111; w[61][65] = 5'b01111; w[61][66] = 5'b01111; w[61][67] = 5'b00000; w[61][68] = 5'b01111; w[61][69] = 5'b01111; w[61][70] = 5'b01111; w[61][71] = 5'b01111; w[61][72] = 5'b00000; w[61][73] = 5'b01111; w[61][74] = 5'b01111; w[61][75] = 5'b01111; w[61][76] = 5'b00000; w[61][77] = 5'b10000; w[61][78] = 5'b01111; w[61][79] = 5'b01111; w[61][80] = 5'b01111; w[61][81] = 5'b00000; w[61][82] = 5'b01111; w[61][83] = 5'b01111; w[61][84] = 5'b01111; w[61][85] = 5'b01111; w[61][86] = 5'b00000; w[61][87] = 5'b01111; w[61][88] = 5'b01111; w[61][89] = 5'b01111; w[61][90] = 5'b00000; w[61][91] = 5'b00000; w[61][92] = 5'b01111; w[61][93] = 5'b01111; w[61][94] = 5'b01111; w[61][95] = 5'b01111; w[61][96] = 5'b01111; w[61][97] = 5'b01111; w[61][98] = 5'b01111; w[61][99] = 5'b01111; w[61][100] = 5'b00000; w[61][101] = 5'b01111; w[61][102] = 5'b01111; w[61][103] = 5'b01111; w[61][104] = 5'b00000; w[61][105] = 5'b00000; w[61][106] = 5'b00000; w[61][107] = 5'b01111; w[61][108] = 5'b01111; w[61][109] = 5'b00000; w[61][110] = 5'b01111; w[61][111] = 5'b01111; w[61][112] = 5'b01111; w[61][113] = 5'b01111; w[61][114] = 5'b00000; w[61][115] = 5'b01111; w[61][116] = 5'b01111; w[61][117] = 5'b01111; w[61][118] = 5'b00000; w[61][119] = 5'b00000; w[61][120] = 5'b01111; w[61][121] = 5'b01111; w[61][122] = 5'b01111; w[61][123] = 5'b00000; w[61][124] = 5'b01111; w[61][125] = 5'b01111; w[61][126] = 5'b01111; w[61][127] = 5'b01111; w[61][128] = 5'b00000; w[61][129] = 5'b01111; w[61][130] = 5'b01111; w[61][131] = 5'b01111; w[61][132] = 5'b10000; w[61][133] = 5'b00000; w[61][134] = 5'b01111; w[61][135] = 5'b01111; w[61][136] = 5'b01111; w[61][137] = 5'b00000; w[61][138] = 5'b01111; w[61][139] = 5'b01111; w[61][140] = 5'b01111; w[61][141] = 5'b01111; w[61][142] = 5'b00000; w[61][143] = 5'b01111; w[61][144] = 5'b01111; w[61][145] = 5'b01111; w[61][146] = 5'b10000; w[61][147] = 5'b00000; w[61][148] = 5'b01111; w[61][149] = 5'b01111; w[61][150] = 5'b01111; w[61][151] = 5'b00000; w[61][152] = 5'b01111; w[61][153] = 5'b01111; w[61][154] = 5'b01111; w[61][155] = 5'b01111; w[61][156] = 5'b01111; w[61][157] = 5'b01111; w[61][158] = 5'b01111; w[61][159] = 5'b10000; w[61][160] = 5'b10000; w[61][161] = 5'b10000; w[61][162] = 5'b00000; w[61][163] = 5'b01111; w[61][164] = 5'b01111; w[61][165] = 5'b01111; w[61][166] = 5'b01111; w[61][167] = 5'b01111; w[61][168] = 5'b01111; w[61][169] = 5'b01111; w[61][170] = 5'b01111; w[61][171] = 5'b01111; w[61][172] = 5'b01111; w[61][173] = 5'b10000; w[61][174] = 5'b10000; w[61][175] = 5'b10000; w[61][176] = 5'b00000; w[61][177] = 5'b01111; w[61][178] = 5'b01111; w[61][179] = 5'b01111; w[61][180] = 5'b01111; w[61][181] = 5'b01111; w[61][182] = 5'b01111; w[61][183] = 5'b01111; w[61][184] = 5'b01111; w[61][185] = 5'b01111; w[61][186] = 5'b01111; w[61][187] = 5'b01111; w[61][188] = 5'b01111; w[61][189] = 5'b01111; w[61][190] = 5'b01111; w[61][191] = 5'b01111; w[61][192] = 5'b01111; w[61][193] = 5'b01111; w[61][194] = 5'b01111; w[61][195] = 5'b01111; w[61][196] = 5'b01111; w[61][197] = 5'b01111; w[61][198] = 5'b01111; w[61][199] = 5'b01111; w[61][200] = 5'b01111; w[61][201] = 5'b01111; w[61][202] = 5'b01111; w[61][203] = 5'b01111; w[61][204] = 5'b01111; w[61][205] = 5'b01111; w[61][206] = 5'b01111; w[61][207] = 5'b01111; w[61][208] = 5'b01111; w[61][209] = 5'b01111; 
w[62][0] = 5'b10000; w[62][1] = 5'b10000; w[62][2] = 5'b10000; w[62][3] = 5'b10000; w[62][4] = 5'b10000; w[62][5] = 5'b10000; w[62][6] = 5'b10000; w[62][7] = 5'b10000; w[62][8] = 5'b10000; w[62][9] = 5'b10000; w[62][10] = 5'b10000; w[62][11] = 5'b10000; w[62][12] = 5'b10000; w[62][13] = 5'b10000; w[62][14] = 5'b10000; w[62][15] = 5'b10000; w[62][16] = 5'b10000; w[62][17] = 5'b10000; w[62][18] = 5'b10000; w[62][19] = 5'b10000; w[62][20] = 5'b10000; w[62][21] = 5'b10000; w[62][22] = 5'b10000; w[62][23] = 5'b10000; w[62][24] = 5'b10000; w[62][25] = 5'b10000; w[62][26] = 5'b10000; w[62][27] = 5'b10000; w[62][28] = 5'b10000; w[62][29] = 5'b10000; w[62][30] = 5'b00000; w[62][31] = 5'b01111; w[62][32] = 5'b00000; w[62][33] = 5'b01111; w[62][34] = 5'b00000; w[62][35] = 5'b00000; w[62][36] = 5'b00000; w[62][37] = 5'b00000; w[62][38] = 5'b01111; w[62][39] = 5'b00000; w[62][40] = 5'b10000; w[62][41] = 5'b10000; w[62][42] = 5'b10000; w[62][43] = 5'b10000; w[62][44] = 5'b00000; w[62][45] = 5'b00000; w[62][46] = 5'b00000; w[62][47] = 5'b01111; w[62][48] = 5'b00000; w[62][49] = 5'b00000; w[62][50] = 5'b00000; w[62][51] = 5'b00000; w[62][52] = 5'b00000; w[62][53] = 5'b00000; w[62][54] = 5'b10000; w[62][55] = 5'b10000; w[62][56] = 5'b10000; w[62][57] = 5'b10000; w[62][58] = 5'b10000; w[62][59] = 5'b10000; w[62][60] = 5'b10000; w[62][61] = 5'b00000; w[62][62] = 5'b00000; w[62][63] = 5'b01111; w[62][64] = 5'b10000; w[62][65] = 5'b10000; w[62][66] = 5'b10000; w[62][67] = 5'b10000; w[62][68] = 5'b10000; w[62][69] = 5'b10000; w[62][70] = 5'b10000; w[62][71] = 5'b10000; w[62][72] = 5'b10000; w[62][73] = 5'b10000; w[62][74] = 5'b00000; w[62][75] = 5'b00000; w[62][76] = 5'b01111; w[62][77] = 5'b01111; w[62][78] = 5'b10000; w[62][79] = 5'b00000; w[62][80] = 5'b10000; w[62][81] = 5'b10000; w[62][82] = 5'b10000; w[62][83] = 5'b10000; w[62][84] = 5'b10000; w[62][85] = 5'b10000; w[62][86] = 5'b10000; w[62][87] = 5'b10000; w[62][88] = 5'b00000; w[62][89] = 5'b00000; w[62][90] = 5'b01111; w[62][91] = 5'b01111; w[62][92] = 5'b10000; w[62][93] = 5'b00000; w[62][94] = 5'b00000; w[62][95] = 5'b10000; w[62][96] = 5'b10000; w[62][97] = 5'b10000; w[62][98] = 5'b10000; w[62][99] = 5'b10000; w[62][100] = 5'b10000; w[62][101] = 5'b10000; w[62][102] = 5'b00000; w[62][103] = 5'b10000; w[62][104] = 5'b01111; w[62][105] = 5'b01111; w[62][106] = 5'b10000; w[62][107] = 5'b10000; w[62][108] = 5'b10000; w[62][109] = 5'b10000; w[62][110] = 5'b10000; w[62][111] = 5'b10000; w[62][112] = 5'b10000; w[62][113] = 5'b10000; w[62][114] = 5'b10000; w[62][115] = 5'b10000; w[62][116] = 5'b00000; w[62][117] = 5'b10000; w[62][118] = 5'b01111; w[62][119] = 5'b01111; w[62][120] = 5'b10000; w[62][121] = 5'b10000; w[62][122] = 5'b10000; w[62][123] = 5'b10000; w[62][124] = 5'b10000; w[62][125] = 5'b10000; w[62][126] = 5'b10000; w[62][127] = 5'b10000; w[62][128] = 5'b10000; w[62][129] = 5'b10000; w[62][130] = 5'b00000; w[62][131] = 5'b10000; w[62][132] = 5'b01111; w[62][133] = 5'b01111; w[62][134] = 5'b00000; w[62][135] = 5'b00000; w[62][136] = 5'b10000; w[62][137] = 5'b10000; w[62][138] = 5'b10000; w[62][139] = 5'b10000; w[62][140] = 5'b10000; w[62][141] = 5'b10000; w[62][142] = 5'b10000; w[62][143] = 5'b10000; w[62][144] = 5'b10000; w[62][145] = 5'b10000; w[62][146] = 5'b01111; w[62][147] = 5'b01111; w[62][148] = 5'b00000; w[62][149] = 5'b10000; w[62][150] = 5'b10000; w[62][151] = 5'b10000; w[62][152] = 5'b10000; w[62][153] = 5'b10000; w[62][154] = 5'b10000; w[62][155] = 5'b10000; w[62][156] = 5'b10000; w[62][157] = 5'b10000; w[62][158] = 5'b10000; w[62][159] = 5'b10000; w[62][160] = 5'b00000; w[62][161] = 5'b00000; w[62][162] = 5'b00000; w[62][163] = 5'b10000; w[62][164] = 5'b10000; w[62][165] = 5'b10000; w[62][166] = 5'b10000; w[62][167] = 5'b10000; w[62][168] = 5'b10000; w[62][169] = 5'b10000; w[62][170] = 5'b10000; w[62][171] = 5'b00000; w[62][172] = 5'b10000; w[62][173] = 5'b10000; w[62][174] = 5'b00000; w[62][175] = 5'b00000; w[62][176] = 5'b00000; w[62][177] = 5'b10000; w[62][178] = 5'b00000; w[62][179] = 5'b10000; w[62][180] = 5'b10000; w[62][181] = 5'b10000; w[62][182] = 5'b10000; w[62][183] = 5'b10000; w[62][184] = 5'b10000; w[62][185] = 5'b10000; w[62][186] = 5'b10000; w[62][187] = 5'b10000; w[62][188] = 5'b10000; w[62][189] = 5'b10000; w[62][190] = 5'b10000; w[62][191] = 5'b10000; w[62][192] = 5'b10000; w[62][193] = 5'b10000; w[62][194] = 5'b10000; w[62][195] = 5'b10000; w[62][196] = 5'b10000; w[62][197] = 5'b10000; w[62][198] = 5'b10000; w[62][199] = 5'b10000; w[62][200] = 5'b10000; w[62][201] = 5'b10000; w[62][202] = 5'b10000; w[62][203] = 5'b10000; w[62][204] = 5'b10000; w[62][205] = 5'b10000; w[62][206] = 5'b10000; w[62][207] = 5'b10000; w[62][208] = 5'b10000; w[62][209] = 5'b10000; 
w[63][0] = 5'b00000; w[63][1] = 5'b00000; w[63][2] = 5'b00000; w[63][3] = 5'b00000; w[63][4] = 5'b00000; w[63][5] = 5'b00000; w[63][6] = 5'b00000; w[63][7] = 5'b00000; w[63][8] = 5'b00000; w[63][9] = 5'b00000; w[63][10] = 5'b00000; w[63][11] = 5'b00000; w[63][12] = 5'b00000; w[63][13] = 5'b00000; w[63][14] = 5'b00000; w[63][15] = 5'b00000; w[63][16] = 5'b00000; w[63][17] = 5'b00000; w[63][18] = 5'b00000; w[63][19] = 5'b00000; w[63][20] = 5'b00000; w[63][21] = 5'b00000; w[63][22] = 5'b00000; w[63][23] = 5'b00000; w[63][24] = 5'b00000; w[63][25] = 5'b00000; w[63][26] = 5'b00000; w[63][27] = 5'b00000; w[63][28] = 5'b00000; w[63][29] = 5'b00000; w[63][30] = 5'b01111; w[63][31] = 5'b00000; w[63][32] = 5'b10000; w[63][33] = 5'b00000; w[63][34] = 5'b01111; w[63][35] = 5'b01111; w[63][36] = 5'b01111; w[63][37] = 5'b10000; w[63][38] = 5'b00000; w[63][39] = 5'b01111; w[63][40] = 5'b00000; w[63][41] = 5'b00000; w[63][42] = 5'b00000; w[63][43] = 5'b00000; w[63][44] = 5'b01111; w[63][45] = 5'b10000; w[63][46] = 5'b10000; w[63][47] = 5'b00000; w[63][48] = 5'b01111; w[63][49] = 5'b01111; w[63][50] = 5'b01111; w[63][51] = 5'b10000; w[63][52] = 5'b10000; w[63][53] = 5'b01111; w[63][54] = 5'b00000; w[63][55] = 5'b00000; w[63][56] = 5'b00000; w[63][57] = 5'b00000; w[63][58] = 5'b10000; w[63][59] = 5'b10000; w[63][60] = 5'b10000; w[63][61] = 5'b10000; w[63][62] = 5'b01111; w[63][63] = 5'b00000; w[63][64] = 5'b00000; w[63][65] = 5'b10000; w[63][66] = 5'b10000; w[63][67] = 5'b10000; w[63][68] = 5'b00000; w[63][69] = 5'b00000; w[63][70] = 5'b00000; w[63][71] = 5'b00000; w[63][72] = 5'b10000; w[63][73] = 5'b10000; w[63][74] = 5'b10000; w[63][75] = 5'b10000; w[63][76] = 5'b01111; w[63][77] = 5'b01111; w[63][78] = 5'b00000; w[63][79] = 5'b10000; w[63][80] = 5'b10000; w[63][81] = 5'b10000; w[63][82] = 5'b00000; w[63][83] = 5'b00000; w[63][84] = 5'b00000; w[63][85] = 5'b00000; w[63][86] = 5'b10000; w[63][87] = 5'b10000; w[63][88] = 5'b10000; w[63][89] = 5'b10000; w[63][90] = 5'b01111; w[63][91] = 5'b01111; w[63][92] = 5'b00000; w[63][93] = 5'b10000; w[63][94] = 5'b10000; w[63][95] = 5'b00000; w[63][96] = 5'b00000; w[63][97] = 5'b00000; w[63][98] = 5'b00000; w[63][99] = 5'b00000; w[63][100] = 5'b10000; w[63][101] = 5'b10000; w[63][102] = 5'b10000; w[63][103] = 5'b00000; w[63][104] = 5'b01111; w[63][105] = 5'b01111; w[63][106] = 5'b10000; w[63][107] = 5'b10000; w[63][108] = 5'b10000; w[63][109] = 5'b10000; w[63][110] = 5'b00000; w[63][111] = 5'b00000; w[63][112] = 5'b00000; w[63][113] = 5'b00000; w[63][114] = 5'b10000; w[63][115] = 5'b10000; w[63][116] = 5'b10000; w[63][117] = 5'b00000; w[63][118] = 5'b01111; w[63][119] = 5'b01111; w[63][120] = 5'b10000; w[63][121] = 5'b10000; w[63][122] = 5'b10000; w[63][123] = 5'b10000; w[63][124] = 5'b00000; w[63][125] = 5'b00000; w[63][126] = 5'b00000; w[63][127] = 5'b00000; w[63][128] = 5'b10000; w[63][129] = 5'b10000; w[63][130] = 5'b10000; w[63][131] = 5'b00000; w[63][132] = 5'b01111; w[63][133] = 5'b01111; w[63][134] = 5'b10000; w[63][135] = 5'b10000; w[63][136] = 5'b10000; w[63][137] = 5'b10000; w[63][138] = 5'b00000; w[63][139] = 5'b00000; w[63][140] = 5'b00000; w[63][141] = 5'b00000; w[63][142] = 5'b10000; w[63][143] = 5'b10000; w[63][144] = 5'b10000; w[63][145] = 5'b00000; w[63][146] = 5'b01111; w[63][147] = 5'b01111; w[63][148] = 5'b10000; w[63][149] = 5'b10000; w[63][150] = 5'b10000; w[63][151] = 5'b10000; w[63][152] = 5'b00000; w[63][153] = 5'b00000; w[63][154] = 5'b00000; w[63][155] = 5'b00000; w[63][156] = 5'b00000; w[63][157] = 5'b10000; w[63][158] = 5'b10000; w[63][159] = 5'b00000; w[63][160] = 5'b01111; w[63][161] = 5'b01111; w[63][162] = 5'b10000; w[63][163] = 5'b10000; w[63][164] = 5'b10000; w[63][165] = 5'b00000; w[63][166] = 5'b00000; w[63][167] = 5'b00000; w[63][168] = 5'b00000; w[63][169] = 5'b00000; w[63][170] = 5'b00000; w[63][171] = 5'b10000; w[63][172] = 5'b10000; w[63][173] = 5'b00000; w[63][174] = 5'b01111; w[63][175] = 5'b01111; w[63][176] = 5'b10000; w[63][177] = 5'b10000; w[63][178] = 5'b10000; w[63][179] = 5'b00000; w[63][180] = 5'b00000; w[63][181] = 5'b00000; w[63][182] = 5'b00000; w[63][183] = 5'b00000; w[63][184] = 5'b00000; w[63][185] = 5'b00000; w[63][186] = 5'b00000; w[63][187] = 5'b00000; w[63][188] = 5'b00000; w[63][189] = 5'b00000; w[63][190] = 5'b00000; w[63][191] = 5'b00000; w[63][192] = 5'b00000; w[63][193] = 5'b00000; w[63][194] = 5'b00000; w[63][195] = 5'b00000; w[63][196] = 5'b00000; w[63][197] = 5'b00000; w[63][198] = 5'b00000; w[63][199] = 5'b00000; w[63][200] = 5'b00000; w[63][201] = 5'b00000; w[63][202] = 5'b00000; w[63][203] = 5'b00000; w[63][204] = 5'b00000; w[63][205] = 5'b00000; w[63][206] = 5'b00000; w[63][207] = 5'b00000; w[63][208] = 5'b00000; w[63][209] = 5'b00000; 
w[64][0] = 5'b01111; w[64][1] = 5'b01111; w[64][2] = 5'b01111; w[64][3] = 5'b01111; w[64][4] = 5'b01111; w[64][5] = 5'b01111; w[64][6] = 5'b01111; w[64][7] = 5'b01111; w[64][8] = 5'b01111; w[64][9] = 5'b01111; w[64][10] = 5'b01111; w[64][11] = 5'b01111; w[64][12] = 5'b01111; w[64][13] = 5'b01111; w[64][14] = 5'b01111; w[64][15] = 5'b01111; w[64][16] = 5'b01111; w[64][17] = 5'b01111; w[64][18] = 5'b01111; w[64][19] = 5'b01111; w[64][20] = 5'b01111; w[64][21] = 5'b01111; w[64][22] = 5'b01111; w[64][23] = 5'b01111; w[64][24] = 5'b01111; w[64][25] = 5'b01111; w[64][26] = 5'b01111; w[64][27] = 5'b01111; w[64][28] = 5'b01111; w[64][29] = 5'b01111; w[64][30] = 5'b01111; w[64][31] = 5'b00000; w[64][32] = 5'b10000; w[64][33] = 5'b10000; w[64][34] = 5'b10000; w[64][35] = 5'b10000; w[64][36] = 5'b10000; w[64][37] = 5'b10000; w[64][38] = 5'b00000; w[64][39] = 5'b01111; w[64][40] = 5'b01111; w[64][41] = 5'b01111; w[64][42] = 5'b01111; w[64][43] = 5'b01111; w[64][44] = 5'b01111; w[64][45] = 5'b10000; w[64][46] = 5'b10000; w[64][47] = 5'b10000; w[64][48] = 5'b10000; w[64][49] = 5'b10000; w[64][50] = 5'b10000; w[64][51] = 5'b10000; w[64][52] = 5'b10000; w[64][53] = 5'b01111; w[64][54] = 5'b01111; w[64][55] = 5'b01111; w[64][56] = 5'b01111; w[64][57] = 5'b01111; w[64][58] = 5'b01111; w[64][59] = 5'b00000; w[64][60] = 5'b00000; w[64][61] = 5'b01111; w[64][62] = 5'b10000; w[64][63] = 5'b00000; w[64][64] = 5'b00000; w[64][65] = 5'b00000; w[64][66] = 5'b00000; w[64][67] = 5'b01111; w[64][68] = 5'b01111; w[64][69] = 5'b01111; w[64][70] = 5'b01111; w[64][71] = 5'b01111; w[64][72] = 5'b01111; w[64][73] = 5'b00000; w[64][74] = 5'b01111; w[64][75] = 5'b01111; w[64][76] = 5'b10000; w[64][77] = 5'b00000; w[64][78] = 5'b01111; w[64][79] = 5'b01111; w[64][80] = 5'b00000; w[64][81] = 5'b01111; w[64][82] = 5'b01111; w[64][83] = 5'b01111; w[64][84] = 5'b01111; w[64][85] = 5'b01111; w[64][86] = 5'b01111; w[64][87] = 5'b00000; w[64][88] = 5'b01111; w[64][89] = 5'b01111; w[64][90] = 5'b10000; w[64][91] = 5'b10000; w[64][92] = 5'b01111; w[64][93] = 5'b01111; w[64][94] = 5'b01111; w[64][95] = 5'b01111; w[64][96] = 5'b01111; w[64][97] = 5'b01111; w[64][98] = 5'b01111; w[64][99] = 5'b01111; w[64][100] = 5'b01111; w[64][101] = 5'b00000; w[64][102] = 5'b01111; w[64][103] = 5'b01111; w[64][104] = 5'b10000; w[64][105] = 5'b10000; w[64][106] = 5'b01111; w[64][107] = 5'b00000; w[64][108] = 5'b00000; w[64][109] = 5'b01111; w[64][110] = 5'b01111; w[64][111] = 5'b01111; w[64][112] = 5'b01111; w[64][113] = 5'b01111; w[64][114] = 5'b01111; w[64][115] = 5'b00000; w[64][116] = 5'b01111; w[64][117] = 5'b01111; w[64][118] = 5'b10000; w[64][119] = 5'b10000; w[64][120] = 5'b00000; w[64][121] = 5'b00000; w[64][122] = 5'b00000; w[64][123] = 5'b01111; w[64][124] = 5'b01111; w[64][125] = 5'b01111; w[64][126] = 5'b01111; w[64][127] = 5'b01111; w[64][128] = 5'b01111; w[64][129] = 5'b00000; w[64][130] = 5'b01111; w[64][131] = 5'b01111; w[64][132] = 5'b00000; w[64][133] = 5'b10000; w[64][134] = 5'b01111; w[64][135] = 5'b01111; w[64][136] = 5'b00000; w[64][137] = 5'b01111; w[64][138] = 5'b01111; w[64][139] = 5'b01111; w[64][140] = 5'b01111; w[64][141] = 5'b01111; w[64][142] = 5'b01111; w[64][143] = 5'b00000; w[64][144] = 5'b00000; w[64][145] = 5'b01111; w[64][146] = 5'b00000; w[64][147] = 5'b10000; w[64][148] = 5'b01111; w[64][149] = 5'b00000; w[64][150] = 5'b00000; w[64][151] = 5'b01111; w[64][152] = 5'b01111; w[64][153] = 5'b01111; w[64][154] = 5'b01111; w[64][155] = 5'b01111; w[64][156] = 5'b01111; w[64][157] = 5'b00000; w[64][158] = 5'b00000; w[64][159] = 5'b00000; w[64][160] = 5'b10000; w[64][161] = 5'b10000; w[64][162] = 5'b10000; w[64][163] = 5'b00000; w[64][164] = 5'b00000; w[64][165] = 5'b01111; w[64][166] = 5'b01111; w[64][167] = 5'b01111; w[64][168] = 5'b01111; w[64][169] = 5'b01111; w[64][170] = 5'b01111; w[64][171] = 5'b01111; w[64][172] = 5'b00000; w[64][173] = 5'b00000; w[64][174] = 5'b10000; w[64][175] = 5'b10000; w[64][176] = 5'b10000; w[64][177] = 5'b00000; w[64][178] = 5'b01111; w[64][179] = 5'b01111; w[64][180] = 5'b01111; w[64][181] = 5'b01111; w[64][182] = 5'b01111; w[64][183] = 5'b01111; w[64][184] = 5'b01111; w[64][185] = 5'b01111; w[64][186] = 5'b01111; w[64][187] = 5'b01111; w[64][188] = 5'b01111; w[64][189] = 5'b01111; w[64][190] = 5'b01111; w[64][191] = 5'b01111; w[64][192] = 5'b01111; w[64][193] = 5'b01111; w[64][194] = 5'b01111; w[64][195] = 5'b01111; w[64][196] = 5'b01111; w[64][197] = 5'b01111; w[64][198] = 5'b01111; w[64][199] = 5'b01111; w[64][200] = 5'b01111; w[64][201] = 5'b01111; w[64][202] = 5'b01111; w[64][203] = 5'b01111; w[64][204] = 5'b01111; w[64][205] = 5'b01111; w[64][206] = 5'b01111; w[64][207] = 5'b01111; w[64][208] = 5'b01111; w[64][209] = 5'b01111; 
w[65][0] = 5'b00000; w[65][1] = 5'b00000; w[65][2] = 5'b00000; w[65][3] = 5'b00000; w[65][4] = 5'b00000; w[65][5] = 5'b00000; w[65][6] = 5'b00000; w[65][7] = 5'b00000; w[65][8] = 5'b00000; w[65][9] = 5'b00000; w[65][10] = 5'b00000; w[65][11] = 5'b00000; w[65][12] = 5'b00000; w[65][13] = 5'b00000; w[65][14] = 5'b00000; w[65][15] = 5'b00000; w[65][16] = 5'b00000; w[65][17] = 5'b00000; w[65][18] = 5'b00000; w[65][19] = 5'b00000; w[65][20] = 5'b00000; w[65][21] = 5'b00000; w[65][22] = 5'b00000; w[65][23] = 5'b00000; w[65][24] = 5'b00000; w[65][25] = 5'b00000; w[65][26] = 5'b00000; w[65][27] = 5'b00000; w[65][28] = 5'b00000; w[65][29] = 5'b00000; w[65][30] = 5'b10000; w[65][31] = 5'b00000; w[65][32] = 5'b01111; w[65][33] = 5'b00000; w[65][34] = 5'b10000; w[65][35] = 5'b10000; w[65][36] = 5'b10000; w[65][37] = 5'b01111; w[65][38] = 5'b00000; w[65][39] = 5'b10000; w[65][40] = 5'b00000; w[65][41] = 5'b00000; w[65][42] = 5'b00000; w[65][43] = 5'b00000; w[65][44] = 5'b10000; w[65][45] = 5'b01111; w[65][46] = 5'b01111; w[65][47] = 5'b00000; w[65][48] = 5'b10000; w[65][49] = 5'b10000; w[65][50] = 5'b10000; w[65][51] = 5'b01111; w[65][52] = 5'b01111; w[65][53] = 5'b10000; w[65][54] = 5'b00000; w[65][55] = 5'b00000; w[65][56] = 5'b00000; w[65][57] = 5'b00000; w[65][58] = 5'b01111; w[65][59] = 5'b01111; w[65][60] = 5'b01111; w[65][61] = 5'b01111; w[65][62] = 5'b10000; w[65][63] = 5'b10000; w[65][64] = 5'b00000; w[65][65] = 5'b00000; w[65][66] = 5'b01111; w[65][67] = 5'b01111; w[65][68] = 5'b00000; w[65][69] = 5'b00000; w[65][70] = 5'b00000; w[65][71] = 5'b00000; w[65][72] = 5'b01111; w[65][73] = 5'b01111; w[65][74] = 5'b01111; w[65][75] = 5'b01111; w[65][76] = 5'b10000; w[65][77] = 5'b10000; w[65][78] = 5'b00000; w[65][79] = 5'b01111; w[65][80] = 5'b01111; w[65][81] = 5'b01111; w[65][82] = 5'b00000; w[65][83] = 5'b00000; w[65][84] = 5'b00000; w[65][85] = 5'b00000; w[65][86] = 5'b01111; w[65][87] = 5'b01111; w[65][88] = 5'b01111; w[65][89] = 5'b01111; w[65][90] = 5'b10000; w[65][91] = 5'b10000; w[65][92] = 5'b00000; w[65][93] = 5'b01111; w[65][94] = 5'b01111; w[65][95] = 5'b00000; w[65][96] = 5'b00000; w[65][97] = 5'b00000; w[65][98] = 5'b00000; w[65][99] = 5'b00000; w[65][100] = 5'b01111; w[65][101] = 5'b01111; w[65][102] = 5'b01111; w[65][103] = 5'b00000; w[65][104] = 5'b10000; w[65][105] = 5'b10000; w[65][106] = 5'b01111; w[65][107] = 5'b01111; w[65][108] = 5'b01111; w[65][109] = 5'b01111; w[65][110] = 5'b00000; w[65][111] = 5'b00000; w[65][112] = 5'b00000; w[65][113] = 5'b00000; w[65][114] = 5'b01111; w[65][115] = 5'b01111; w[65][116] = 5'b01111; w[65][117] = 5'b00000; w[65][118] = 5'b10000; w[65][119] = 5'b10000; w[65][120] = 5'b01111; w[65][121] = 5'b01111; w[65][122] = 5'b01111; w[65][123] = 5'b01111; w[65][124] = 5'b00000; w[65][125] = 5'b00000; w[65][126] = 5'b00000; w[65][127] = 5'b00000; w[65][128] = 5'b01111; w[65][129] = 5'b01111; w[65][130] = 5'b01111; w[65][131] = 5'b00000; w[65][132] = 5'b10000; w[65][133] = 5'b10000; w[65][134] = 5'b01111; w[65][135] = 5'b01111; w[65][136] = 5'b01111; w[65][137] = 5'b01111; w[65][138] = 5'b00000; w[65][139] = 5'b00000; w[65][140] = 5'b00000; w[65][141] = 5'b00000; w[65][142] = 5'b01111; w[65][143] = 5'b01111; w[65][144] = 5'b01111; w[65][145] = 5'b00000; w[65][146] = 5'b10000; w[65][147] = 5'b10000; w[65][148] = 5'b01111; w[65][149] = 5'b01111; w[65][150] = 5'b01111; w[65][151] = 5'b01111; w[65][152] = 5'b00000; w[65][153] = 5'b00000; w[65][154] = 5'b00000; w[65][155] = 5'b00000; w[65][156] = 5'b00000; w[65][157] = 5'b01111; w[65][158] = 5'b01111; w[65][159] = 5'b00000; w[65][160] = 5'b10000; w[65][161] = 5'b10000; w[65][162] = 5'b01111; w[65][163] = 5'b01111; w[65][164] = 5'b01111; w[65][165] = 5'b00000; w[65][166] = 5'b00000; w[65][167] = 5'b00000; w[65][168] = 5'b00000; w[65][169] = 5'b00000; w[65][170] = 5'b00000; w[65][171] = 5'b01111; w[65][172] = 5'b01111; w[65][173] = 5'b00000; w[65][174] = 5'b10000; w[65][175] = 5'b10000; w[65][176] = 5'b01111; w[65][177] = 5'b01111; w[65][178] = 5'b01111; w[65][179] = 5'b00000; w[65][180] = 5'b00000; w[65][181] = 5'b00000; w[65][182] = 5'b00000; w[65][183] = 5'b00000; w[65][184] = 5'b00000; w[65][185] = 5'b00000; w[65][186] = 5'b00000; w[65][187] = 5'b00000; w[65][188] = 5'b00000; w[65][189] = 5'b00000; w[65][190] = 5'b00000; w[65][191] = 5'b00000; w[65][192] = 5'b00000; w[65][193] = 5'b00000; w[65][194] = 5'b00000; w[65][195] = 5'b00000; w[65][196] = 5'b00000; w[65][197] = 5'b00000; w[65][198] = 5'b00000; w[65][199] = 5'b00000; w[65][200] = 5'b00000; w[65][201] = 5'b00000; w[65][202] = 5'b00000; w[65][203] = 5'b00000; w[65][204] = 5'b00000; w[65][205] = 5'b00000; w[65][206] = 5'b00000; w[65][207] = 5'b00000; w[65][208] = 5'b00000; w[65][209] = 5'b00000; 
w[66][0] = 5'b00000; w[66][1] = 5'b00000; w[66][2] = 5'b00000; w[66][3] = 5'b00000; w[66][4] = 5'b00000; w[66][5] = 5'b00000; w[66][6] = 5'b00000; w[66][7] = 5'b00000; w[66][8] = 5'b00000; w[66][9] = 5'b00000; w[66][10] = 5'b00000; w[66][11] = 5'b00000; w[66][12] = 5'b00000; w[66][13] = 5'b00000; w[66][14] = 5'b00000; w[66][15] = 5'b00000; w[66][16] = 5'b00000; w[66][17] = 5'b00000; w[66][18] = 5'b00000; w[66][19] = 5'b00000; w[66][20] = 5'b00000; w[66][21] = 5'b00000; w[66][22] = 5'b00000; w[66][23] = 5'b00000; w[66][24] = 5'b00000; w[66][25] = 5'b00000; w[66][26] = 5'b00000; w[66][27] = 5'b00000; w[66][28] = 5'b00000; w[66][29] = 5'b00000; w[66][30] = 5'b10000; w[66][31] = 5'b00000; w[66][32] = 5'b01111; w[66][33] = 5'b00000; w[66][34] = 5'b10000; w[66][35] = 5'b10000; w[66][36] = 5'b10000; w[66][37] = 5'b01111; w[66][38] = 5'b00000; w[66][39] = 5'b10000; w[66][40] = 5'b00000; w[66][41] = 5'b00000; w[66][42] = 5'b00000; w[66][43] = 5'b00000; w[66][44] = 5'b10000; w[66][45] = 5'b01111; w[66][46] = 5'b01111; w[66][47] = 5'b00000; w[66][48] = 5'b10000; w[66][49] = 5'b10000; w[66][50] = 5'b10000; w[66][51] = 5'b01111; w[66][52] = 5'b01111; w[66][53] = 5'b10000; w[66][54] = 5'b00000; w[66][55] = 5'b00000; w[66][56] = 5'b00000; w[66][57] = 5'b00000; w[66][58] = 5'b01111; w[66][59] = 5'b01111; w[66][60] = 5'b01111; w[66][61] = 5'b01111; w[66][62] = 5'b10000; w[66][63] = 5'b10000; w[66][64] = 5'b00000; w[66][65] = 5'b01111; w[66][66] = 5'b00000; w[66][67] = 5'b01111; w[66][68] = 5'b00000; w[66][69] = 5'b00000; w[66][70] = 5'b00000; w[66][71] = 5'b00000; w[66][72] = 5'b01111; w[66][73] = 5'b01111; w[66][74] = 5'b01111; w[66][75] = 5'b01111; w[66][76] = 5'b10000; w[66][77] = 5'b10000; w[66][78] = 5'b00000; w[66][79] = 5'b01111; w[66][80] = 5'b01111; w[66][81] = 5'b01111; w[66][82] = 5'b00000; w[66][83] = 5'b00000; w[66][84] = 5'b00000; w[66][85] = 5'b00000; w[66][86] = 5'b01111; w[66][87] = 5'b01111; w[66][88] = 5'b01111; w[66][89] = 5'b01111; w[66][90] = 5'b10000; w[66][91] = 5'b10000; w[66][92] = 5'b00000; w[66][93] = 5'b01111; w[66][94] = 5'b01111; w[66][95] = 5'b00000; w[66][96] = 5'b00000; w[66][97] = 5'b00000; w[66][98] = 5'b00000; w[66][99] = 5'b00000; w[66][100] = 5'b01111; w[66][101] = 5'b01111; w[66][102] = 5'b01111; w[66][103] = 5'b00000; w[66][104] = 5'b10000; w[66][105] = 5'b10000; w[66][106] = 5'b01111; w[66][107] = 5'b01111; w[66][108] = 5'b01111; w[66][109] = 5'b01111; w[66][110] = 5'b00000; w[66][111] = 5'b00000; w[66][112] = 5'b00000; w[66][113] = 5'b00000; w[66][114] = 5'b01111; w[66][115] = 5'b01111; w[66][116] = 5'b01111; w[66][117] = 5'b00000; w[66][118] = 5'b10000; w[66][119] = 5'b10000; w[66][120] = 5'b01111; w[66][121] = 5'b01111; w[66][122] = 5'b01111; w[66][123] = 5'b01111; w[66][124] = 5'b00000; w[66][125] = 5'b00000; w[66][126] = 5'b00000; w[66][127] = 5'b00000; w[66][128] = 5'b01111; w[66][129] = 5'b01111; w[66][130] = 5'b01111; w[66][131] = 5'b00000; w[66][132] = 5'b10000; w[66][133] = 5'b10000; w[66][134] = 5'b01111; w[66][135] = 5'b01111; w[66][136] = 5'b01111; w[66][137] = 5'b01111; w[66][138] = 5'b00000; w[66][139] = 5'b00000; w[66][140] = 5'b00000; w[66][141] = 5'b00000; w[66][142] = 5'b01111; w[66][143] = 5'b01111; w[66][144] = 5'b01111; w[66][145] = 5'b00000; w[66][146] = 5'b10000; w[66][147] = 5'b10000; w[66][148] = 5'b01111; w[66][149] = 5'b01111; w[66][150] = 5'b01111; w[66][151] = 5'b01111; w[66][152] = 5'b00000; w[66][153] = 5'b00000; w[66][154] = 5'b00000; w[66][155] = 5'b00000; w[66][156] = 5'b00000; w[66][157] = 5'b01111; w[66][158] = 5'b01111; w[66][159] = 5'b00000; w[66][160] = 5'b10000; w[66][161] = 5'b10000; w[66][162] = 5'b01111; w[66][163] = 5'b01111; w[66][164] = 5'b01111; w[66][165] = 5'b00000; w[66][166] = 5'b00000; w[66][167] = 5'b00000; w[66][168] = 5'b00000; w[66][169] = 5'b00000; w[66][170] = 5'b00000; w[66][171] = 5'b01111; w[66][172] = 5'b01111; w[66][173] = 5'b00000; w[66][174] = 5'b10000; w[66][175] = 5'b10000; w[66][176] = 5'b01111; w[66][177] = 5'b01111; w[66][178] = 5'b01111; w[66][179] = 5'b00000; w[66][180] = 5'b00000; w[66][181] = 5'b00000; w[66][182] = 5'b00000; w[66][183] = 5'b00000; w[66][184] = 5'b00000; w[66][185] = 5'b00000; w[66][186] = 5'b00000; w[66][187] = 5'b00000; w[66][188] = 5'b00000; w[66][189] = 5'b00000; w[66][190] = 5'b00000; w[66][191] = 5'b00000; w[66][192] = 5'b00000; w[66][193] = 5'b00000; w[66][194] = 5'b00000; w[66][195] = 5'b00000; w[66][196] = 5'b00000; w[66][197] = 5'b00000; w[66][198] = 5'b00000; w[66][199] = 5'b00000; w[66][200] = 5'b00000; w[66][201] = 5'b00000; w[66][202] = 5'b00000; w[66][203] = 5'b00000; w[66][204] = 5'b00000; w[66][205] = 5'b00000; w[66][206] = 5'b00000; w[66][207] = 5'b00000; w[66][208] = 5'b00000; w[66][209] = 5'b00000; 
w[67][0] = 5'b01111; w[67][1] = 5'b01111; w[67][2] = 5'b01111; w[67][3] = 5'b01111; w[67][4] = 5'b01111; w[67][5] = 5'b01111; w[67][6] = 5'b01111; w[67][7] = 5'b01111; w[67][8] = 5'b01111; w[67][9] = 5'b01111; w[67][10] = 5'b01111; w[67][11] = 5'b01111; w[67][12] = 5'b01111; w[67][13] = 5'b01111; w[67][14] = 5'b01111; w[67][15] = 5'b01111; w[67][16] = 5'b01111; w[67][17] = 5'b01111; w[67][18] = 5'b01111; w[67][19] = 5'b01111; w[67][20] = 5'b01111; w[67][21] = 5'b01111; w[67][22] = 5'b01111; w[67][23] = 5'b01111; w[67][24] = 5'b01111; w[67][25] = 5'b01111; w[67][26] = 5'b01111; w[67][27] = 5'b01111; w[67][28] = 5'b01111; w[67][29] = 5'b01111; w[67][30] = 5'b00000; w[67][31] = 5'b10000; w[67][32] = 5'b00000; w[67][33] = 5'b10000; w[67][34] = 5'b00000; w[67][35] = 5'b00000; w[67][36] = 5'b00000; w[67][37] = 5'b00000; w[67][38] = 5'b10000; w[67][39] = 5'b00000; w[67][40] = 5'b01111; w[67][41] = 5'b01111; w[67][42] = 5'b01111; w[67][43] = 5'b01111; w[67][44] = 5'b00000; w[67][45] = 5'b00000; w[67][46] = 5'b00000; w[67][47] = 5'b10000; w[67][48] = 5'b00000; w[67][49] = 5'b00000; w[67][50] = 5'b00000; w[67][51] = 5'b00000; w[67][52] = 5'b00000; w[67][53] = 5'b00000; w[67][54] = 5'b01111; w[67][55] = 5'b01111; w[67][56] = 5'b01111; w[67][57] = 5'b01111; w[67][58] = 5'b01111; w[67][59] = 5'b01111; w[67][60] = 5'b01111; w[67][61] = 5'b00000; w[67][62] = 5'b10000; w[67][63] = 5'b10000; w[67][64] = 5'b01111; w[67][65] = 5'b01111; w[67][66] = 5'b01111; w[67][67] = 5'b00000; w[67][68] = 5'b01111; w[67][69] = 5'b01111; w[67][70] = 5'b01111; w[67][71] = 5'b01111; w[67][72] = 5'b01111; w[67][73] = 5'b01111; w[67][74] = 5'b00000; w[67][75] = 5'b00000; w[67][76] = 5'b10000; w[67][77] = 5'b10000; w[67][78] = 5'b01111; w[67][79] = 5'b00000; w[67][80] = 5'b01111; w[67][81] = 5'b01111; w[67][82] = 5'b01111; w[67][83] = 5'b01111; w[67][84] = 5'b01111; w[67][85] = 5'b01111; w[67][86] = 5'b01111; w[67][87] = 5'b01111; w[67][88] = 5'b00000; w[67][89] = 5'b00000; w[67][90] = 5'b10000; w[67][91] = 5'b10000; w[67][92] = 5'b01111; w[67][93] = 5'b00000; w[67][94] = 5'b00000; w[67][95] = 5'b01111; w[67][96] = 5'b01111; w[67][97] = 5'b01111; w[67][98] = 5'b01111; w[67][99] = 5'b01111; w[67][100] = 5'b01111; w[67][101] = 5'b01111; w[67][102] = 5'b00000; w[67][103] = 5'b01111; w[67][104] = 5'b10000; w[67][105] = 5'b10000; w[67][106] = 5'b01111; w[67][107] = 5'b01111; w[67][108] = 5'b01111; w[67][109] = 5'b01111; w[67][110] = 5'b01111; w[67][111] = 5'b01111; w[67][112] = 5'b01111; w[67][113] = 5'b01111; w[67][114] = 5'b01111; w[67][115] = 5'b01111; w[67][116] = 5'b00000; w[67][117] = 5'b01111; w[67][118] = 5'b10000; w[67][119] = 5'b10000; w[67][120] = 5'b01111; w[67][121] = 5'b01111; w[67][122] = 5'b01111; w[67][123] = 5'b01111; w[67][124] = 5'b01111; w[67][125] = 5'b01111; w[67][126] = 5'b01111; w[67][127] = 5'b01111; w[67][128] = 5'b01111; w[67][129] = 5'b01111; w[67][130] = 5'b00000; w[67][131] = 5'b01111; w[67][132] = 5'b10000; w[67][133] = 5'b10000; w[67][134] = 5'b00000; w[67][135] = 5'b00000; w[67][136] = 5'b01111; w[67][137] = 5'b01111; w[67][138] = 5'b01111; w[67][139] = 5'b01111; w[67][140] = 5'b01111; w[67][141] = 5'b01111; w[67][142] = 5'b01111; w[67][143] = 5'b01111; w[67][144] = 5'b01111; w[67][145] = 5'b01111; w[67][146] = 5'b10000; w[67][147] = 5'b10000; w[67][148] = 5'b00000; w[67][149] = 5'b01111; w[67][150] = 5'b01111; w[67][151] = 5'b01111; w[67][152] = 5'b01111; w[67][153] = 5'b01111; w[67][154] = 5'b01111; w[67][155] = 5'b01111; w[67][156] = 5'b01111; w[67][157] = 5'b01111; w[67][158] = 5'b01111; w[67][159] = 5'b01111; w[67][160] = 5'b00000; w[67][161] = 5'b00000; w[67][162] = 5'b00000; w[67][163] = 5'b01111; w[67][164] = 5'b01111; w[67][165] = 5'b01111; w[67][166] = 5'b01111; w[67][167] = 5'b01111; w[67][168] = 5'b01111; w[67][169] = 5'b01111; w[67][170] = 5'b01111; w[67][171] = 5'b00000; w[67][172] = 5'b01111; w[67][173] = 5'b01111; w[67][174] = 5'b00000; w[67][175] = 5'b00000; w[67][176] = 5'b00000; w[67][177] = 5'b01111; w[67][178] = 5'b00000; w[67][179] = 5'b01111; w[67][180] = 5'b01111; w[67][181] = 5'b01111; w[67][182] = 5'b01111; w[67][183] = 5'b01111; w[67][184] = 5'b01111; w[67][185] = 5'b01111; w[67][186] = 5'b01111; w[67][187] = 5'b01111; w[67][188] = 5'b01111; w[67][189] = 5'b01111; w[67][190] = 5'b01111; w[67][191] = 5'b01111; w[67][192] = 5'b01111; w[67][193] = 5'b01111; w[67][194] = 5'b01111; w[67][195] = 5'b01111; w[67][196] = 5'b01111; w[67][197] = 5'b01111; w[67][198] = 5'b01111; w[67][199] = 5'b01111; w[67][200] = 5'b01111; w[67][201] = 5'b01111; w[67][202] = 5'b01111; w[67][203] = 5'b01111; w[67][204] = 5'b01111; w[67][205] = 5'b01111; w[67][206] = 5'b01111; w[67][207] = 5'b01111; w[67][208] = 5'b01111; w[67][209] = 5'b01111; 
w[68][0] = 5'b01111; w[68][1] = 5'b01111; w[68][2] = 5'b01111; w[68][3] = 5'b01111; w[68][4] = 5'b01111; w[68][5] = 5'b01111; w[68][6] = 5'b01111; w[68][7] = 5'b01111; w[68][8] = 5'b01111; w[68][9] = 5'b01111; w[68][10] = 5'b01111; w[68][11] = 5'b01111; w[68][12] = 5'b01111; w[68][13] = 5'b01111; w[68][14] = 5'b01111; w[68][15] = 5'b01111; w[68][16] = 5'b01111; w[68][17] = 5'b01111; w[68][18] = 5'b01111; w[68][19] = 5'b01111; w[68][20] = 5'b01111; w[68][21] = 5'b01111; w[68][22] = 5'b01111; w[68][23] = 5'b01111; w[68][24] = 5'b01111; w[68][25] = 5'b01111; w[68][26] = 5'b01111; w[68][27] = 5'b01111; w[68][28] = 5'b01111; w[68][29] = 5'b01111; w[68][30] = 5'b01111; w[68][31] = 5'b00000; w[68][32] = 5'b10000; w[68][33] = 5'b10000; w[68][34] = 5'b10000; w[68][35] = 5'b10000; w[68][36] = 5'b10000; w[68][37] = 5'b10000; w[68][38] = 5'b00000; w[68][39] = 5'b01111; w[68][40] = 5'b01111; w[68][41] = 5'b01111; w[68][42] = 5'b01111; w[68][43] = 5'b01111; w[68][44] = 5'b01111; w[68][45] = 5'b10000; w[68][46] = 5'b10000; w[68][47] = 5'b10000; w[68][48] = 5'b10000; w[68][49] = 5'b10000; w[68][50] = 5'b10000; w[68][51] = 5'b10000; w[68][52] = 5'b10000; w[68][53] = 5'b01111; w[68][54] = 5'b01111; w[68][55] = 5'b01111; w[68][56] = 5'b01111; w[68][57] = 5'b01111; w[68][58] = 5'b01111; w[68][59] = 5'b00000; w[68][60] = 5'b00000; w[68][61] = 5'b01111; w[68][62] = 5'b10000; w[68][63] = 5'b00000; w[68][64] = 5'b01111; w[68][65] = 5'b00000; w[68][66] = 5'b00000; w[68][67] = 5'b01111; w[68][68] = 5'b00000; w[68][69] = 5'b01111; w[68][70] = 5'b01111; w[68][71] = 5'b01111; w[68][72] = 5'b01111; w[68][73] = 5'b00000; w[68][74] = 5'b01111; w[68][75] = 5'b01111; w[68][76] = 5'b10000; w[68][77] = 5'b00000; w[68][78] = 5'b01111; w[68][79] = 5'b01111; w[68][80] = 5'b00000; w[68][81] = 5'b01111; w[68][82] = 5'b01111; w[68][83] = 5'b01111; w[68][84] = 5'b01111; w[68][85] = 5'b01111; w[68][86] = 5'b01111; w[68][87] = 5'b00000; w[68][88] = 5'b01111; w[68][89] = 5'b01111; w[68][90] = 5'b10000; w[68][91] = 5'b10000; w[68][92] = 5'b01111; w[68][93] = 5'b01111; w[68][94] = 5'b01111; w[68][95] = 5'b01111; w[68][96] = 5'b01111; w[68][97] = 5'b01111; w[68][98] = 5'b01111; w[68][99] = 5'b01111; w[68][100] = 5'b01111; w[68][101] = 5'b00000; w[68][102] = 5'b01111; w[68][103] = 5'b01111; w[68][104] = 5'b10000; w[68][105] = 5'b10000; w[68][106] = 5'b01111; w[68][107] = 5'b00000; w[68][108] = 5'b00000; w[68][109] = 5'b01111; w[68][110] = 5'b01111; w[68][111] = 5'b01111; w[68][112] = 5'b01111; w[68][113] = 5'b01111; w[68][114] = 5'b01111; w[68][115] = 5'b00000; w[68][116] = 5'b01111; w[68][117] = 5'b01111; w[68][118] = 5'b10000; w[68][119] = 5'b10000; w[68][120] = 5'b00000; w[68][121] = 5'b00000; w[68][122] = 5'b00000; w[68][123] = 5'b01111; w[68][124] = 5'b01111; w[68][125] = 5'b01111; w[68][126] = 5'b01111; w[68][127] = 5'b01111; w[68][128] = 5'b01111; w[68][129] = 5'b00000; w[68][130] = 5'b01111; w[68][131] = 5'b01111; w[68][132] = 5'b00000; w[68][133] = 5'b10000; w[68][134] = 5'b01111; w[68][135] = 5'b01111; w[68][136] = 5'b00000; w[68][137] = 5'b01111; w[68][138] = 5'b01111; w[68][139] = 5'b01111; w[68][140] = 5'b01111; w[68][141] = 5'b01111; w[68][142] = 5'b01111; w[68][143] = 5'b00000; w[68][144] = 5'b00000; w[68][145] = 5'b01111; w[68][146] = 5'b00000; w[68][147] = 5'b10000; w[68][148] = 5'b01111; w[68][149] = 5'b00000; w[68][150] = 5'b00000; w[68][151] = 5'b01111; w[68][152] = 5'b01111; w[68][153] = 5'b01111; w[68][154] = 5'b01111; w[68][155] = 5'b01111; w[68][156] = 5'b01111; w[68][157] = 5'b00000; w[68][158] = 5'b00000; w[68][159] = 5'b00000; w[68][160] = 5'b10000; w[68][161] = 5'b10000; w[68][162] = 5'b10000; w[68][163] = 5'b00000; w[68][164] = 5'b00000; w[68][165] = 5'b01111; w[68][166] = 5'b01111; w[68][167] = 5'b01111; w[68][168] = 5'b01111; w[68][169] = 5'b01111; w[68][170] = 5'b01111; w[68][171] = 5'b01111; w[68][172] = 5'b00000; w[68][173] = 5'b00000; w[68][174] = 5'b10000; w[68][175] = 5'b10000; w[68][176] = 5'b10000; w[68][177] = 5'b00000; w[68][178] = 5'b01111; w[68][179] = 5'b01111; w[68][180] = 5'b01111; w[68][181] = 5'b01111; w[68][182] = 5'b01111; w[68][183] = 5'b01111; w[68][184] = 5'b01111; w[68][185] = 5'b01111; w[68][186] = 5'b01111; w[68][187] = 5'b01111; w[68][188] = 5'b01111; w[68][189] = 5'b01111; w[68][190] = 5'b01111; w[68][191] = 5'b01111; w[68][192] = 5'b01111; w[68][193] = 5'b01111; w[68][194] = 5'b01111; w[68][195] = 5'b01111; w[68][196] = 5'b01111; w[68][197] = 5'b01111; w[68][198] = 5'b01111; w[68][199] = 5'b01111; w[68][200] = 5'b01111; w[68][201] = 5'b01111; w[68][202] = 5'b01111; w[68][203] = 5'b01111; w[68][204] = 5'b01111; w[68][205] = 5'b01111; w[68][206] = 5'b01111; w[68][207] = 5'b01111; w[68][208] = 5'b01111; w[68][209] = 5'b01111; 
w[69][0] = 5'b01111; w[69][1] = 5'b01111; w[69][2] = 5'b01111; w[69][3] = 5'b01111; w[69][4] = 5'b01111; w[69][5] = 5'b01111; w[69][6] = 5'b01111; w[69][7] = 5'b01111; w[69][8] = 5'b01111; w[69][9] = 5'b01111; w[69][10] = 5'b01111; w[69][11] = 5'b01111; w[69][12] = 5'b01111; w[69][13] = 5'b01111; w[69][14] = 5'b01111; w[69][15] = 5'b01111; w[69][16] = 5'b01111; w[69][17] = 5'b01111; w[69][18] = 5'b01111; w[69][19] = 5'b01111; w[69][20] = 5'b01111; w[69][21] = 5'b01111; w[69][22] = 5'b01111; w[69][23] = 5'b01111; w[69][24] = 5'b01111; w[69][25] = 5'b01111; w[69][26] = 5'b01111; w[69][27] = 5'b01111; w[69][28] = 5'b01111; w[69][29] = 5'b01111; w[69][30] = 5'b01111; w[69][31] = 5'b00000; w[69][32] = 5'b10000; w[69][33] = 5'b10000; w[69][34] = 5'b10000; w[69][35] = 5'b10000; w[69][36] = 5'b10000; w[69][37] = 5'b10000; w[69][38] = 5'b00000; w[69][39] = 5'b01111; w[69][40] = 5'b01111; w[69][41] = 5'b01111; w[69][42] = 5'b01111; w[69][43] = 5'b01111; w[69][44] = 5'b01111; w[69][45] = 5'b10000; w[69][46] = 5'b10000; w[69][47] = 5'b10000; w[69][48] = 5'b10000; w[69][49] = 5'b10000; w[69][50] = 5'b10000; w[69][51] = 5'b10000; w[69][52] = 5'b10000; w[69][53] = 5'b01111; w[69][54] = 5'b01111; w[69][55] = 5'b01111; w[69][56] = 5'b01111; w[69][57] = 5'b01111; w[69][58] = 5'b01111; w[69][59] = 5'b00000; w[69][60] = 5'b00000; w[69][61] = 5'b01111; w[69][62] = 5'b10000; w[69][63] = 5'b00000; w[69][64] = 5'b01111; w[69][65] = 5'b00000; w[69][66] = 5'b00000; w[69][67] = 5'b01111; w[69][68] = 5'b01111; w[69][69] = 5'b00000; w[69][70] = 5'b01111; w[69][71] = 5'b01111; w[69][72] = 5'b01111; w[69][73] = 5'b00000; w[69][74] = 5'b01111; w[69][75] = 5'b01111; w[69][76] = 5'b10000; w[69][77] = 5'b00000; w[69][78] = 5'b01111; w[69][79] = 5'b01111; w[69][80] = 5'b00000; w[69][81] = 5'b01111; w[69][82] = 5'b01111; w[69][83] = 5'b01111; w[69][84] = 5'b01111; w[69][85] = 5'b01111; w[69][86] = 5'b01111; w[69][87] = 5'b00000; w[69][88] = 5'b01111; w[69][89] = 5'b01111; w[69][90] = 5'b10000; w[69][91] = 5'b10000; w[69][92] = 5'b01111; w[69][93] = 5'b01111; w[69][94] = 5'b01111; w[69][95] = 5'b01111; w[69][96] = 5'b01111; w[69][97] = 5'b01111; w[69][98] = 5'b01111; w[69][99] = 5'b01111; w[69][100] = 5'b01111; w[69][101] = 5'b00000; w[69][102] = 5'b01111; w[69][103] = 5'b01111; w[69][104] = 5'b10000; w[69][105] = 5'b10000; w[69][106] = 5'b01111; w[69][107] = 5'b00000; w[69][108] = 5'b00000; w[69][109] = 5'b01111; w[69][110] = 5'b01111; w[69][111] = 5'b01111; w[69][112] = 5'b01111; w[69][113] = 5'b01111; w[69][114] = 5'b01111; w[69][115] = 5'b00000; w[69][116] = 5'b01111; w[69][117] = 5'b01111; w[69][118] = 5'b10000; w[69][119] = 5'b10000; w[69][120] = 5'b00000; w[69][121] = 5'b00000; w[69][122] = 5'b00000; w[69][123] = 5'b01111; w[69][124] = 5'b01111; w[69][125] = 5'b01111; w[69][126] = 5'b01111; w[69][127] = 5'b01111; w[69][128] = 5'b01111; w[69][129] = 5'b00000; w[69][130] = 5'b01111; w[69][131] = 5'b01111; w[69][132] = 5'b00000; w[69][133] = 5'b10000; w[69][134] = 5'b01111; w[69][135] = 5'b01111; w[69][136] = 5'b00000; w[69][137] = 5'b01111; w[69][138] = 5'b01111; w[69][139] = 5'b01111; w[69][140] = 5'b01111; w[69][141] = 5'b01111; w[69][142] = 5'b01111; w[69][143] = 5'b00000; w[69][144] = 5'b00000; w[69][145] = 5'b01111; w[69][146] = 5'b00000; w[69][147] = 5'b10000; w[69][148] = 5'b01111; w[69][149] = 5'b00000; w[69][150] = 5'b00000; w[69][151] = 5'b01111; w[69][152] = 5'b01111; w[69][153] = 5'b01111; w[69][154] = 5'b01111; w[69][155] = 5'b01111; w[69][156] = 5'b01111; w[69][157] = 5'b00000; w[69][158] = 5'b00000; w[69][159] = 5'b00000; w[69][160] = 5'b10000; w[69][161] = 5'b10000; w[69][162] = 5'b10000; w[69][163] = 5'b00000; w[69][164] = 5'b00000; w[69][165] = 5'b01111; w[69][166] = 5'b01111; w[69][167] = 5'b01111; w[69][168] = 5'b01111; w[69][169] = 5'b01111; w[69][170] = 5'b01111; w[69][171] = 5'b01111; w[69][172] = 5'b00000; w[69][173] = 5'b00000; w[69][174] = 5'b10000; w[69][175] = 5'b10000; w[69][176] = 5'b10000; w[69][177] = 5'b00000; w[69][178] = 5'b01111; w[69][179] = 5'b01111; w[69][180] = 5'b01111; w[69][181] = 5'b01111; w[69][182] = 5'b01111; w[69][183] = 5'b01111; w[69][184] = 5'b01111; w[69][185] = 5'b01111; w[69][186] = 5'b01111; w[69][187] = 5'b01111; w[69][188] = 5'b01111; w[69][189] = 5'b01111; w[69][190] = 5'b01111; w[69][191] = 5'b01111; w[69][192] = 5'b01111; w[69][193] = 5'b01111; w[69][194] = 5'b01111; w[69][195] = 5'b01111; w[69][196] = 5'b01111; w[69][197] = 5'b01111; w[69][198] = 5'b01111; w[69][199] = 5'b01111; w[69][200] = 5'b01111; w[69][201] = 5'b01111; w[69][202] = 5'b01111; w[69][203] = 5'b01111; w[69][204] = 5'b01111; w[69][205] = 5'b01111; w[69][206] = 5'b01111; w[69][207] = 5'b01111; w[69][208] = 5'b01111; w[69][209] = 5'b01111; 
w[70][0] = 5'b01111; w[70][1] = 5'b01111; w[70][2] = 5'b01111; w[70][3] = 5'b01111; w[70][4] = 5'b01111; w[70][5] = 5'b01111; w[70][6] = 5'b01111; w[70][7] = 5'b01111; w[70][8] = 5'b01111; w[70][9] = 5'b01111; w[70][10] = 5'b01111; w[70][11] = 5'b01111; w[70][12] = 5'b01111; w[70][13] = 5'b01111; w[70][14] = 5'b01111; w[70][15] = 5'b01111; w[70][16] = 5'b01111; w[70][17] = 5'b01111; w[70][18] = 5'b01111; w[70][19] = 5'b01111; w[70][20] = 5'b01111; w[70][21] = 5'b01111; w[70][22] = 5'b01111; w[70][23] = 5'b01111; w[70][24] = 5'b01111; w[70][25] = 5'b01111; w[70][26] = 5'b01111; w[70][27] = 5'b01111; w[70][28] = 5'b01111; w[70][29] = 5'b01111; w[70][30] = 5'b01111; w[70][31] = 5'b00000; w[70][32] = 5'b10000; w[70][33] = 5'b10000; w[70][34] = 5'b10000; w[70][35] = 5'b10000; w[70][36] = 5'b10000; w[70][37] = 5'b10000; w[70][38] = 5'b00000; w[70][39] = 5'b01111; w[70][40] = 5'b01111; w[70][41] = 5'b01111; w[70][42] = 5'b01111; w[70][43] = 5'b01111; w[70][44] = 5'b01111; w[70][45] = 5'b10000; w[70][46] = 5'b10000; w[70][47] = 5'b10000; w[70][48] = 5'b10000; w[70][49] = 5'b10000; w[70][50] = 5'b10000; w[70][51] = 5'b10000; w[70][52] = 5'b10000; w[70][53] = 5'b01111; w[70][54] = 5'b01111; w[70][55] = 5'b01111; w[70][56] = 5'b01111; w[70][57] = 5'b01111; w[70][58] = 5'b01111; w[70][59] = 5'b00000; w[70][60] = 5'b00000; w[70][61] = 5'b01111; w[70][62] = 5'b10000; w[70][63] = 5'b00000; w[70][64] = 5'b01111; w[70][65] = 5'b00000; w[70][66] = 5'b00000; w[70][67] = 5'b01111; w[70][68] = 5'b01111; w[70][69] = 5'b01111; w[70][70] = 5'b00000; w[70][71] = 5'b01111; w[70][72] = 5'b01111; w[70][73] = 5'b00000; w[70][74] = 5'b01111; w[70][75] = 5'b01111; w[70][76] = 5'b10000; w[70][77] = 5'b00000; w[70][78] = 5'b01111; w[70][79] = 5'b01111; w[70][80] = 5'b00000; w[70][81] = 5'b01111; w[70][82] = 5'b01111; w[70][83] = 5'b01111; w[70][84] = 5'b01111; w[70][85] = 5'b01111; w[70][86] = 5'b01111; w[70][87] = 5'b00000; w[70][88] = 5'b01111; w[70][89] = 5'b01111; w[70][90] = 5'b10000; w[70][91] = 5'b10000; w[70][92] = 5'b01111; w[70][93] = 5'b01111; w[70][94] = 5'b01111; w[70][95] = 5'b01111; w[70][96] = 5'b01111; w[70][97] = 5'b01111; w[70][98] = 5'b01111; w[70][99] = 5'b01111; w[70][100] = 5'b01111; w[70][101] = 5'b00000; w[70][102] = 5'b01111; w[70][103] = 5'b01111; w[70][104] = 5'b10000; w[70][105] = 5'b10000; w[70][106] = 5'b01111; w[70][107] = 5'b00000; w[70][108] = 5'b00000; w[70][109] = 5'b01111; w[70][110] = 5'b01111; w[70][111] = 5'b01111; w[70][112] = 5'b01111; w[70][113] = 5'b01111; w[70][114] = 5'b01111; w[70][115] = 5'b00000; w[70][116] = 5'b01111; w[70][117] = 5'b01111; w[70][118] = 5'b10000; w[70][119] = 5'b10000; w[70][120] = 5'b00000; w[70][121] = 5'b00000; w[70][122] = 5'b00000; w[70][123] = 5'b01111; w[70][124] = 5'b01111; w[70][125] = 5'b01111; w[70][126] = 5'b01111; w[70][127] = 5'b01111; w[70][128] = 5'b01111; w[70][129] = 5'b00000; w[70][130] = 5'b01111; w[70][131] = 5'b01111; w[70][132] = 5'b00000; w[70][133] = 5'b10000; w[70][134] = 5'b01111; w[70][135] = 5'b01111; w[70][136] = 5'b00000; w[70][137] = 5'b01111; w[70][138] = 5'b01111; w[70][139] = 5'b01111; w[70][140] = 5'b01111; w[70][141] = 5'b01111; w[70][142] = 5'b01111; w[70][143] = 5'b00000; w[70][144] = 5'b00000; w[70][145] = 5'b01111; w[70][146] = 5'b00000; w[70][147] = 5'b10000; w[70][148] = 5'b01111; w[70][149] = 5'b00000; w[70][150] = 5'b00000; w[70][151] = 5'b01111; w[70][152] = 5'b01111; w[70][153] = 5'b01111; w[70][154] = 5'b01111; w[70][155] = 5'b01111; w[70][156] = 5'b01111; w[70][157] = 5'b00000; w[70][158] = 5'b00000; w[70][159] = 5'b00000; w[70][160] = 5'b10000; w[70][161] = 5'b10000; w[70][162] = 5'b10000; w[70][163] = 5'b00000; w[70][164] = 5'b00000; w[70][165] = 5'b01111; w[70][166] = 5'b01111; w[70][167] = 5'b01111; w[70][168] = 5'b01111; w[70][169] = 5'b01111; w[70][170] = 5'b01111; w[70][171] = 5'b01111; w[70][172] = 5'b00000; w[70][173] = 5'b00000; w[70][174] = 5'b10000; w[70][175] = 5'b10000; w[70][176] = 5'b10000; w[70][177] = 5'b00000; w[70][178] = 5'b01111; w[70][179] = 5'b01111; w[70][180] = 5'b01111; w[70][181] = 5'b01111; w[70][182] = 5'b01111; w[70][183] = 5'b01111; w[70][184] = 5'b01111; w[70][185] = 5'b01111; w[70][186] = 5'b01111; w[70][187] = 5'b01111; w[70][188] = 5'b01111; w[70][189] = 5'b01111; w[70][190] = 5'b01111; w[70][191] = 5'b01111; w[70][192] = 5'b01111; w[70][193] = 5'b01111; w[70][194] = 5'b01111; w[70][195] = 5'b01111; w[70][196] = 5'b01111; w[70][197] = 5'b01111; w[70][198] = 5'b01111; w[70][199] = 5'b01111; w[70][200] = 5'b01111; w[70][201] = 5'b01111; w[70][202] = 5'b01111; w[70][203] = 5'b01111; w[70][204] = 5'b01111; w[70][205] = 5'b01111; w[70][206] = 5'b01111; w[70][207] = 5'b01111; w[70][208] = 5'b01111; w[70][209] = 5'b01111; 
w[71][0] = 5'b01111; w[71][1] = 5'b01111; w[71][2] = 5'b01111; w[71][3] = 5'b01111; w[71][4] = 5'b01111; w[71][5] = 5'b01111; w[71][6] = 5'b01111; w[71][7] = 5'b01111; w[71][8] = 5'b01111; w[71][9] = 5'b01111; w[71][10] = 5'b01111; w[71][11] = 5'b01111; w[71][12] = 5'b01111; w[71][13] = 5'b01111; w[71][14] = 5'b01111; w[71][15] = 5'b01111; w[71][16] = 5'b01111; w[71][17] = 5'b01111; w[71][18] = 5'b01111; w[71][19] = 5'b01111; w[71][20] = 5'b01111; w[71][21] = 5'b01111; w[71][22] = 5'b01111; w[71][23] = 5'b01111; w[71][24] = 5'b01111; w[71][25] = 5'b01111; w[71][26] = 5'b01111; w[71][27] = 5'b01111; w[71][28] = 5'b01111; w[71][29] = 5'b01111; w[71][30] = 5'b01111; w[71][31] = 5'b00000; w[71][32] = 5'b10000; w[71][33] = 5'b10000; w[71][34] = 5'b10000; w[71][35] = 5'b10000; w[71][36] = 5'b10000; w[71][37] = 5'b10000; w[71][38] = 5'b00000; w[71][39] = 5'b01111; w[71][40] = 5'b01111; w[71][41] = 5'b01111; w[71][42] = 5'b01111; w[71][43] = 5'b01111; w[71][44] = 5'b01111; w[71][45] = 5'b10000; w[71][46] = 5'b10000; w[71][47] = 5'b10000; w[71][48] = 5'b10000; w[71][49] = 5'b10000; w[71][50] = 5'b10000; w[71][51] = 5'b10000; w[71][52] = 5'b10000; w[71][53] = 5'b01111; w[71][54] = 5'b01111; w[71][55] = 5'b01111; w[71][56] = 5'b01111; w[71][57] = 5'b01111; w[71][58] = 5'b01111; w[71][59] = 5'b00000; w[71][60] = 5'b00000; w[71][61] = 5'b01111; w[71][62] = 5'b10000; w[71][63] = 5'b00000; w[71][64] = 5'b01111; w[71][65] = 5'b00000; w[71][66] = 5'b00000; w[71][67] = 5'b01111; w[71][68] = 5'b01111; w[71][69] = 5'b01111; w[71][70] = 5'b01111; w[71][71] = 5'b00000; w[71][72] = 5'b01111; w[71][73] = 5'b00000; w[71][74] = 5'b01111; w[71][75] = 5'b01111; w[71][76] = 5'b10000; w[71][77] = 5'b00000; w[71][78] = 5'b01111; w[71][79] = 5'b01111; w[71][80] = 5'b00000; w[71][81] = 5'b01111; w[71][82] = 5'b01111; w[71][83] = 5'b01111; w[71][84] = 5'b01111; w[71][85] = 5'b01111; w[71][86] = 5'b01111; w[71][87] = 5'b00000; w[71][88] = 5'b01111; w[71][89] = 5'b01111; w[71][90] = 5'b10000; w[71][91] = 5'b10000; w[71][92] = 5'b01111; w[71][93] = 5'b01111; w[71][94] = 5'b01111; w[71][95] = 5'b01111; w[71][96] = 5'b01111; w[71][97] = 5'b01111; w[71][98] = 5'b01111; w[71][99] = 5'b01111; w[71][100] = 5'b01111; w[71][101] = 5'b00000; w[71][102] = 5'b01111; w[71][103] = 5'b01111; w[71][104] = 5'b10000; w[71][105] = 5'b10000; w[71][106] = 5'b01111; w[71][107] = 5'b00000; w[71][108] = 5'b00000; w[71][109] = 5'b01111; w[71][110] = 5'b01111; w[71][111] = 5'b01111; w[71][112] = 5'b01111; w[71][113] = 5'b01111; w[71][114] = 5'b01111; w[71][115] = 5'b00000; w[71][116] = 5'b01111; w[71][117] = 5'b01111; w[71][118] = 5'b10000; w[71][119] = 5'b10000; w[71][120] = 5'b00000; w[71][121] = 5'b00000; w[71][122] = 5'b00000; w[71][123] = 5'b01111; w[71][124] = 5'b01111; w[71][125] = 5'b01111; w[71][126] = 5'b01111; w[71][127] = 5'b01111; w[71][128] = 5'b01111; w[71][129] = 5'b00000; w[71][130] = 5'b01111; w[71][131] = 5'b01111; w[71][132] = 5'b00000; w[71][133] = 5'b10000; w[71][134] = 5'b01111; w[71][135] = 5'b01111; w[71][136] = 5'b00000; w[71][137] = 5'b01111; w[71][138] = 5'b01111; w[71][139] = 5'b01111; w[71][140] = 5'b01111; w[71][141] = 5'b01111; w[71][142] = 5'b01111; w[71][143] = 5'b00000; w[71][144] = 5'b00000; w[71][145] = 5'b01111; w[71][146] = 5'b00000; w[71][147] = 5'b10000; w[71][148] = 5'b01111; w[71][149] = 5'b00000; w[71][150] = 5'b00000; w[71][151] = 5'b01111; w[71][152] = 5'b01111; w[71][153] = 5'b01111; w[71][154] = 5'b01111; w[71][155] = 5'b01111; w[71][156] = 5'b01111; w[71][157] = 5'b00000; w[71][158] = 5'b00000; w[71][159] = 5'b00000; w[71][160] = 5'b10000; w[71][161] = 5'b10000; w[71][162] = 5'b10000; w[71][163] = 5'b00000; w[71][164] = 5'b00000; w[71][165] = 5'b01111; w[71][166] = 5'b01111; w[71][167] = 5'b01111; w[71][168] = 5'b01111; w[71][169] = 5'b01111; w[71][170] = 5'b01111; w[71][171] = 5'b01111; w[71][172] = 5'b00000; w[71][173] = 5'b00000; w[71][174] = 5'b10000; w[71][175] = 5'b10000; w[71][176] = 5'b10000; w[71][177] = 5'b00000; w[71][178] = 5'b01111; w[71][179] = 5'b01111; w[71][180] = 5'b01111; w[71][181] = 5'b01111; w[71][182] = 5'b01111; w[71][183] = 5'b01111; w[71][184] = 5'b01111; w[71][185] = 5'b01111; w[71][186] = 5'b01111; w[71][187] = 5'b01111; w[71][188] = 5'b01111; w[71][189] = 5'b01111; w[71][190] = 5'b01111; w[71][191] = 5'b01111; w[71][192] = 5'b01111; w[71][193] = 5'b01111; w[71][194] = 5'b01111; w[71][195] = 5'b01111; w[71][196] = 5'b01111; w[71][197] = 5'b01111; w[71][198] = 5'b01111; w[71][199] = 5'b01111; w[71][200] = 5'b01111; w[71][201] = 5'b01111; w[71][202] = 5'b01111; w[71][203] = 5'b01111; w[71][204] = 5'b01111; w[71][205] = 5'b01111; w[71][206] = 5'b01111; w[71][207] = 5'b01111; w[71][208] = 5'b01111; w[71][209] = 5'b01111; 
w[72][0] = 5'b01111; w[72][1] = 5'b01111; w[72][2] = 5'b01111; w[72][3] = 5'b01111; w[72][4] = 5'b01111; w[72][5] = 5'b01111; w[72][6] = 5'b01111; w[72][7] = 5'b01111; w[72][8] = 5'b01111; w[72][9] = 5'b01111; w[72][10] = 5'b01111; w[72][11] = 5'b01111; w[72][12] = 5'b01111; w[72][13] = 5'b01111; w[72][14] = 5'b01111; w[72][15] = 5'b01111; w[72][16] = 5'b01111; w[72][17] = 5'b01111; w[72][18] = 5'b01111; w[72][19] = 5'b01111; w[72][20] = 5'b01111; w[72][21] = 5'b01111; w[72][22] = 5'b01111; w[72][23] = 5'b01111; w[72][24] = 5'b01111; w[72][25] = 5'b01111; w[72][26] = 5'b01111; w[72][27] = 5'b01111; w[72][28] = 5'b01111; w[72][29] = 5'b01111; w[72][30] = 5'b00000; w[72][31] = 5'b10000; w[72][32] = 5'b00000; w[72][33] = 5'b10000; w[72][34] = 5'b00000; w[72][35] = 5'b00000; w[72][36] = 5'b00000; w[72][37] = 5'b00000; w[72][38] = 5'b10000; w[72][39] = 5'b00000; w[72][40] = 5'b01111; w[72][41] = 5'b01111; w[72][42] = 5'b01111; w[72][43] = 5'b01111; w[72][44] = 5'b00000; w[72][45] = 5'b00000; w[72][46] = 5'b00000; w[72][47] = 5'b10000; w[72][48] = 5'b00000; w[72][49] = 5'b00000; w[72][50] = 5'b00000; w[72][51] = 5'b00000; w[72][52] = 5'b00000; w[72][53] = 5'b00000; w[72][54] = 5'b01111; w[72][55] = 5'b01111; w[72][56] = 5'b01111; w[72][57] = 5'b01111; w[72][58] = 5'b01111; w[72][59] = 5'b01111; w[72][60] = 5'b01111; w[72][61] = 5'b00000; w[72][62] = 5'b10000; w[72][63] = 5'b10000; w[72][64] = 5'b01111; w[72][65] = 5'b01111; w[72][66] = 5'b01111; w[72][67] = 5'b01111; w[72][68] = 5'b01111; w[72][69] = 5'b01111; w[72][70] = 5'b01111; w[72][71] = 5'b01111; w[72][72] = 5'b00000; w[72][73] = 5'b01111; w[72][74] = 5'b00000; w[72][75] = 5'b00000; w[72][76] = 5'b10000; w[72][77] = 5'b10000; w[72][78] = 5'b01111; w[72][79] = 5'b00000; w[72][80] = 5'b01111; w[72][81] = 5'b01111; w[72][82] = 5'b01111; w[72][83] = 5'b01111; w[72][84] = 5'b01111; w[72][85] = 5'b01111; w[72][86] = 5'b01111; w[72][87] = 5'b01111; w[72][88] = 5'b00000; w[72][89] = 5'b00000; w[72][90] = 5'b10000; w[72][91] = 5'b10000; w[72][92] = 5'b01111; w[72][93] = 5'b00000; w[72][94] = 5'b00000; w[72][95] = 5'b01111; w[72][96] = 5'b01111; w[72][97] = 5'b01111; w[72][98] = 5'b01111; w[72][99] = 5'b01111; w[72][100] = 5'b01111; w[72][101] = 5'b01111; w[72][102] = 5'b00000; w[72][103] = 5'b01111; w[72][104] = 5'b10000; w[72][105] = 5'b10000; w[72][106] = 5'b01111; w[72][107] = 5'b01111; w[72][108] = 5'b01111; w[72][109] = 5'b01111; w[72][110] = 5'b01111; w[72][111] = 5'b01111; w[72][112] = 5'b01111; w[72][113] = 5'b01111; w[72][114] = 5'b01111; w[72][115] = 5'b01111; w[72][116] = 5'b00000; w[72][117] = 5'b01111; w[72][118] = 5'b10000; w[72][119] = 5'b10000; w[72][120] = 5'b01111; w[72][121] = 5'b01111; w[72][122] = 5'b01111; w[72][123] = 5'b01111; w[72][124] = 5'b01111; w[72][125] = 5'b01111; w[72][126] = 5'b01111; w[72][127] = 5'b01111; w[72][128] = 5'b01111; w[72][129] = 5'b01111; w[72][130] = 5'b00000; w[72][131] = 5'b01111; w[72][132] = 5'b10000; w[72][133] = 5'b10000; w[72][134] = 5'b00000; w[72][135] = 5'b00000; w[72][136] = 5'b01111; w[72][137] = 5'b01111; w[72][138] = 5'b01111; w[72][139] = 5'b01111; w[72][140] = 5'b01111; w[72][141] = 5'b01111; w[72][142] = 5'b01111; w[72][143] = 5'b01111; w[72][144] = 5'b01111; w[72][145] = 5'b01111; w[72][146] = 5'b10000; w[72][147] = 5'b10000; w[72][148] = 5'b00000; w[72][149] = 5'b01111; w[72][150] = 5'b01111; w[72][151] = 5'b01111; w[72][152] = 5'b01111; w[72][153] = 5'b01111; w[72][154] = 5'b01111; w[72][155] = 5'b01111; w[72][156] = 5'b01111; w[72][157] = 5'b01111; w[72][158] = 5'b01111; w[72][159] = 5'b01111; w[72][160] = 5'b00000; w[72][161] = 5'b00000; w[72][162] = 5'b00000; w[72][163] = 5'b01111; w[72][164] = 5'b01111; w[72][165] = 5'b01111; w[72][166] = 5'b01111; w[72][167] = 5'b01111; w[72][168] = 5'b01111; w[72][169] = 5'b01111; w[72][170] = 5'b01111; w[72][171] = 5'b00000; w[72][172] = 5'b01111; w[72][173] = 5'b01111; w[72][174] = 5'b00000; w[72][175] = 5'b00000; w[72][176] = 5'b00000; w[72][177] = 5'b01111; w[72][178] = 5'b00000; w[72][179] = 5'b01111; w[72][180] = 5'b01111; w[72][181] = 5'b01111; w[72][182] = 5'b01111; w[72][183] = 5'b01111; w[72][184] = 5'b01111; w[72][185] = 5'b01111; w[72][186] = 5'b01111; w[72][187] = 5'b01111; w[72][188] = 5'b01111; w[72][189] = 5'b01111; w[72][190] = 5'b01111; w[72][191] = 5'b01111; w[72][192] = 5'b01111; w[72][193] = 5'b01111; w[72][194] = 5'b01111; w[72][195] = 5'b01111; w[72][196] = 5'b01111; w[72][197] = 5'b01111; w[72][198] = 5'b01111; w[72][199] = 5'b01111; w[72][200] = 5'b01111; w[72][201] = 5'b01111; w[72][202] = 5'b01111; w[72][203] = 5'b01111; w[72][204] = 5'b01111; w[72][205] = 5'b01111; w[72][206] = 5'b01111; w[72][207] = 5'b01111; w[72][208] = 5'b01111; w[72][209] = 5'b01111; 
w[73][0] = 5'b00000; w[73][1] = 5'b00000; w[73][2] = 5'b00000; w[73][3] = 5'b00000; w[73][4] = 5'b00000; w[73][5] = 5'b00000; w[73][6] = 5'b00000; w[73][7] = 5'b00000; w[73][8] = 5'b00000; w[73][9] = 5'b00000; w[73][10] = 5'b00000; w[73][11] = 5'b00000; w[73][12] = 5'b00000; w[73][13] = 5'b00000; w[73][14] = 5'b00000; w[73][15] = 5'b00000; w[73][16] = 5'b00000; w[73][17] = 5'b00000; w[73][18] = 5'b00000; w[73][19] = 5'b00000; w[73][20] = 5'b00000; w[73][21] = 5'b00000; w[73][22] = 5'b00000; w[73][23] = 5'b00000; w[73][24] = 5'b00000; w[73][25] = 5'b00000; w[73][26] = 5'b00000; w[73][27] = 5'b00000; w[73][28] = 5'b00000; w[73][29] = 5'b00000; w[73][30] = 5'b10000; w[73][31] = 5'b00000; w[73][32] = 5'b01111; w[73][33] = 5'b00000; w[73][34] = 5'b10000; w[73][35] = 5'b10000; w[73][36] = 5'b10000; w[73][37] = 5'b01111; w[73][38] = 5'b00000; w[73][39] = 5'b10000; w[73][40] = 5'b00000; w[73][41] = 5'b00000; w[73][42] = 5'b00000; w[73][43] = 5'b00000; w[73][44] = 5'b10000; w[73][45] = 5'b01111; w[73][46] = 5'b01111; w[73][47] = 5'b00000; w[73][48] = 5'b10000; w[73][49] = 5'b10000; w[73][50] = 5'b10000; w[73][51] = 5'b01111; w[73][52] = 5'b01111; w[73][53] = 5'b10000; w[73][54] = 5'b00000; w[73][55] = 5'b00000; w[73][56] = 5'b00000; w[73][57] = 5'b00000; w[73][58] = 5'b01111; w[73][59] = 5'b01111; w[73][60] = 5'b01111; w[73][61] = 5'b01111; w[73][62] = 5'b10000; w[73][63] = 5'b10000; w[73][64] = 5'b00000; w[73][65] = 5'b01111; w[73][66] = 5'b01111; w[73][67] = 5'b01111; w[73][68] = 5'b00000; w[73][69] = 5'b00000; w[73][70] = 5'b00000; w[73][71] = 5'b00000; w[73][72] = 5'b01111; w[73][73] = 5'b00000; w[73][74] = 5'b01111; w[73][75] = 5'b01111; w[73][76] = 5'b10000; w[73][77] = 5'b10000; w[73][78] = 5'b00000; w[73][79] = 5'b01111; w[73][80] = 5'b01111; w[73][81] = 5'b01111; w[73][82] = 5'b00000; w[73][83] = 5'b00000; w[73][84] = 5'b00000; w[73][85] = 5'b00000; w[73][86] = 5'b01111; w[73][87] = 5'b01111; w[73][88] = 5'b01111; w[73][89] = 5'b01111; w[73][90] = 5'b10000; w[73][91] = 5'b10000; w[73][92] = 5'b00000; w[73][93] = 5'b01111; w[73][94] = 5'b01111; w[73][95] = 5'b00000; w[73][96] = 5'b00000; w[73][97] = 5'b00000; w[73][98] = 5'b00000; w[73][99] = 5'b00000; w[73][100] = 5'b01111; w[73][101] = 5'b01111; w[73][102] = 5'b01111; w[73][103] = 5'b00000; w[73][104] = 5'b10000; w[73][105] = 5'b10000; w[73][106] = 5'b01111; w[73][107] = 5'b01111; w[73][108] = 5'b01111; w[73][109] = 5'b01111; w[73][110] = 5'b00000; w[73][111] = 5'b00000; w[73][112] = 5'b00000; w[73][113] = 5'b00000; w[73][114] = 5'b01111; w[73][115] = 5'b01111; w[73][116] = 5'b01111; w[73][117] = 5'b00000; w[73][118] = 5'b10000; w[73][119] = 5'b10000; w[73][120] = 5'b01111; w[73][121] = 5'b01111; w[73][122] = 5'b01111; w[73][123] = 5'b01111; w[73][124] = 5'b00000; w[73][125] = 5'b00000; w[73][126] = 5'b00000; w[73][127] = 5'b00000; w[73][128] = 5'b01111; w[73][129] = 5'b01111; w[73][130] = 5'b01111; w[73][131] = 5'b00000; w[73][132] = 5'b10000; w[73][133] = 5'b10000; w[73][134] = 5'b01111; w[73][135] = 5'b01111; w[73][136] = 5'b01111; w[73][137] = 5'b01111; w[73][138] = 5'b00000; w[73][139] = 5'b00000; w[73][140] = 5'b00000; w[73][141] = 5'b00000; w[73][142] = 5'b01111; w[73][143] = 5'b01111; w[73][144] = 5'b01111; w[73][145] = 5'b00000; w[73][146] = 5'b10000; w[73][147] = 5'b10000; w[73][148] = 5'b01111; w[73][149] = 5'b01111; w[73][150] = 5'b01111; w[73][151] = 5'b01111; w[73][152] = 5'b00000; w[73][153] = 5'b00000; w[73][154] = 5'b00000; w[73][155] = 5'b00000; w[73][156] = 5'b00000; w[73][157] = 5'b01111; w[73][158] = 5'b01111; w[73][159] = 5'b00000; w[73][160] = 5'b10000; w[73][161] = 5'b10000; w[73][162] = 5'b01111; w[73][163] = 5'b01111; w[73][164] = 5'b01111; w[73][165] = 5'b00000; w[73][166] = 5'b00000; w[73][167] = 5'b00000; w[73][168] = 5'b00000; w[73][169] = 5'b00000; w[73][170] = 5'b00000; w[73][171] = 5'b01111; w[73][172] = 5'b01111; w[73][173] = 5'b00000; w[73][174] = 5'b10000; w[73][175] = 5'b10000; w[73][176] = 5'b01111; w[73][177] = 5'b01111; w[73][178] = 5'b01111; w[73][179] = 5'b00000; w[73][180] = 5'b00000; w[73][181] = 5'b00000; w[73][182] = 5'b00000; w[73][183] = 5'b00000; w[73][184] = 5'b00000; w[73][185] = 5'b00000; w[73][186] = 5'b00000; w[73][187] = 5'b00000; w[73][188] = 5'b00000; w[73][189] = 5'b00000; w[73][190] = 5'b00000; w[73][191] = 5'b00000; w[73][192] = 5'b00000; w[73][193] = 5'b00000; w[73][194] = 5'b00000; w[73][195] = 5'b00000; w[73][196] = 5'b00000; w[73][197] = 5'b00000; w[73][198] = 5'b00000; w[73][199] = 5'b00000; w[73][200] = 5'b00000; w[73][201] = 5'b00000; w[73][202] = 5'b00000; w[73][203] = 5'b00000; w[73][204] = 5'b00000; w[73][205] = 5'b00000; w[73][206] = 5'b00000; w[73][207] = 5'b00000; w[73][208] = 5'b00000; w[73][209] = 5'b00000; 
w[74][0] = 5'b01111; w[74][1] = 5'b01111; w[74][2] = 5'b01111; w[74][3] = 5'b01111; w[74][4] = 5'b01111; w[74][5] = 5'b01111; w[74][6] = 5'b01111; w[74][7] = 5'b01111; w[74][8] = 5'b01111; w[74][9] = 5'b01111; w[74][10] = 5'b01111; w[74][11] = 5'b01111; w[74][12] = 5'b01111; w[74][13] = 5'b01111; w[74][14] = 5'b01111; w[74][15] = 5'b01111; w[74][16] = 5'b01111; w[74][17] = 5'b01111; w[74][18] = 5'b01111; w[74][19] = 5'b01111; w[74][20] = 5'b01111; w[74][21] = 5'b01111; w[74][22] = 5'b01111; w[74][23] = 5'b01111; w[74][24] = 5'b01111; w[74][25] = 5'b01111; w[74][26] = 5'b01111; w[74][27] = 5'b01111; w[74][28] = 5'b01111; w[74][29] = 5'b01111; w[74][30] = 5'b00000; w[74][31] = 5'b01111; w[74][32] = 5'b00000; w[74][33] = 5'b10000; w[74][34] = 5'b10000; w[74][35] = 5'b10000; w[74][36] = 5'b10000; w[74][37] = 5'b00000; w[74][38] = 5'b01111; w[74][39] = 5'b00000; w[74][40] = 5'b01111; w[74][41] = 5'b01111; w[74][42] = 5'b01111; w[74][43] = 5'b01111; w[74][44] = 5'b00000; w[74][45] = 5'b00000; w[74][46] = 5'b00000; w[74][47] = 5'b10000; w[74][48] = 5'b10000; w[74][49] = 5'b10000; w[74][50] = 5'b10000; w[74][51] = 5'b00000; w[74][52] = 5'b00000; w[74][53] = 5'b00000; w[74][54] = 5'b01111; w[74][55] = 5'b01111; w[74][56] = 5'b01111; w[74][57] = 5'b01111; w[74][58] = 5'b00000; w[74][59] = 5'b01111; w[74][60] = 5'b01111; w[74][61] = 5'b01111; w[74][62] = 5'b00000; w[74][63] = 5'b10000; w[74][64] = 5'b01111; w[74][65] = 5'b01111; w[74][66] = 5'b01111; w[74][67] = 5'b00000; w[74][68] = 5'b01111; w[74][69] = 5'b01111; w[74][70] = 5'b01111; w[74][71] = 5'b01111; w[74][72] = 5'b00000; w[74][73] = 5'b01111; w[74][74] = 5'b00000; w[74][75] = 5'b01111; w[74][76] = 5'b00000; w[74][77] = 5'b10000; w[74][78] = 5'b01111; w[74][79] = 5'b01111; w[74][80] = 5'b01111; w[74][81] = 5'b00000; w[74][82] = 5'b01111; w[74][83] = 5'b01111; w[74][84] = 5'b01111; w[74][85] = 5'b01111; w[74][86] = 5'b00000; w[74][87] = 5'b01111; w[74][88] = 5'b01111; w[74][89] = 5'b01111; w[74][90] = 5'b00000; w[74][91] = 5'b00000; w[74][92] = 5'b01111; w[74][93] = 5'b01111; w[74][94] = 5'b01111; w[74][95] = 5'b01111; w[74][96] = 5'b01111; w[74][97] = 5'b01111; w[74][98] = 5'b01111; w[74][99] = 5'b01111; w[74][100] = 5'b00000; w[74][101] = 5'b01111; w[74][102] = 5'b01111; w[74][103] = 5'b01111; w[74][104] = 5'b00000; w[74][105] = 5'b00000; w[74][106] = 5'b00000; w[74][107] = 5'b01111; w[74][108] = 5'b01111; w[74][109] = 5'b00000; w[74][110] = 5'b01111; w[74][111] = 5'b01111; w[74][112] = 5'b01111; w[74][113] = 5'b01111; w[74][114] = 5'b00000; w[74][115] = 5'b01111; w[74][116] = 5'b01111; w[74][117] = 5'b01111; w[74][118] = 5'b00000; w[74][119] = 5'b00000; w[74][120] = 5'b01111; w[74][121] = 5'b01111; w[74][122] = 5'b01111; w[74][123] = 5'b00000; w[74][124] = 5'b01111; w[74][125] = 5'b01111; w[74][126] = 5'b01111; w[74][127] = 5'b01111; w[74][128] = 5'b00000; w[74][129] = 5'b01111; w[74][130] = 5'b01111; w[74][131] = 5'b01111; w[74][132] = 5'b10000; w[74][133] = 5'b00000; w[74][134] = 5'b01111; w[74][135] = 5'b01111; w[74][136] = 5'b01111; w[74][137] = 5'b00000; w[74][138] = 5'b01111; w[74][139] = 5'b01111; w[74][140] = 5'b01111; w[74][141] = 5'b01111; w[74][142] = 5'b00000; w[74][143] = 5'b01111; w[74][144] = 5'b01111; w[74][145] = 5'b01111; w[74][146] = 5'b10000; w[74][147] = 5'b00000; w[74][148] = 5'b01111; w[74][149] = 5'b01111; w[74][150] = 5'b01111; w[74][151] = 5'b00000; w[74][152] = 5'b01111; w[74][153] = 5'b01111; w[74][154] = 5'b01111; w[74][155] = 5'b01111; w[74][156] = 5'b01111; w[74][157] = 5'b01111; w[74][158] = 5'b01111; w[74][159] = 5'b10000; w[74][160] = 5'b10000; w[74][161] = 5'b10000; w[74][162] = 5'b00000; w[74][163] = 5'b01111; w[74][164] = 5'b01111; w[74][165] = 5'b01111; w[74][166] = 5'b01111; w[74][167] = 5'b01111; w[74][168] = 5'b01111; w[74][169] = 5'b01111; w[74][170] = 5'b01111; w[74][171] = 5'b01111; w[74][172] = 5'b01111; w[74][173] = 5'b10000; w[74][174] = 5'b10000; w[74][175] = 5'b10000; w[74][176] = 5'b00000; w[74][177] = 5'b01111; w[74][178] = 5'b01111; w[74][179] = 5'b01111; w[74][180] = 5'b01111; w[74][181] = 5'b01111; w[74][182] = 5'b01111; w[74][183] = 5'b01111; w[74][184] = 5'b01111; w[74][185] = 5'b01111; w[74][186] = 5'b01111; w[74][187] = 5'b01111; w[74][188] = 5'b01111; w[74][189] = 5'b01111; w[74][190] = 5'b01111; w[74][191] = 5'b01111; w[74][192] = 5'b01111; w[74][193] = 5'b01111; w[74][194] = 5'b01111; w[74][195] = 5'b01111; w[74][196] = 5'b01111; w[74][197] = 5'b01111; w[74][198] = 5'b01111; w[74][199] = 5'b01111; w[74][200] = 5'b01111; w[74][201] = 5'b01111; w[74][202] = 5'b01111; w[74][203] = 5'b01111; w[74][204] = 5'b01111; w[74][205] = 5'b01111; w[74][206] = 5'b01111; w[74][207] = 5'b01111; w[74][208] = 5'b01111; w[74][209] = 5'b01111; 
w[75][0] = 5'b01111; w[75][1] = 5'b01111; w[75][2] = 5'b01111; w[75][3] = 5'b01111; w[75][4] = 5'b01111; w[75][5] = 5'b01111; w[75][6] = 5'b01111; w[75][7] = 5'b01111; w[75][8] = 5'b01111; w[75][9] = 5'b01111; w[75][10] = 5'b01111; w[75][11] = 5'b01111; w[75][12] = 5'b01111; w[75][13] = 5'b01111; w[75][14] = 5'b01111; w[75][15] = 5'b01111; w[75][16] = 5'b01111; w[75][17] = 5'b01111; w[75][18] = 5'b01111; w[75][19] = 5'b01111; w[75][20] = 5'b01111; w[75][21] = 5'b01111; w[75][22] = 5'b01111; w[75][23] = 5'b01111; w[75][24] = 5'b01111; w[75][25] = 5'b01111; w[75][26] = 5'b01111; w[75][27] = 5'b01111; w[75][28] = 5'b01111; w[75][29] = 5'b01111; w[75][30] = 5'b00000; w[75][31] = 5'b01111; w[75][32] = 5'b00000; w[75][33] = 5'b10000; w[75][34] = 5'b10000; w[75][35] = 5'b10000; w[75][36] = 5'b10000; w[75][37] = 5'b00000; w[75][38] = 5'b01111; w[75][39] = 5'b00000; w[75][40] = 5'b01111; w[75][41] = 5'b01111; w[75][42] = 5'b01111; w[75][43] = 5'b01111; w[75][44] = 5'b00000; w[75][45] = 5'b00000; w[75][46] = 5'b00000; w[75][47] = 5'b10000; w[75][48] = 5'b10000; w[75][49] = 5'b10000; w[75][50] = 5'b10000; w[75][51] = 5'b00000; w[75][52] = 5'b00000; w[75][53] = 5'b00000; w[75][54] = 5'b01111; w[75][55] = 5'b01111; w[75][56] = 5'b01111; w[75][57] = 5'b01111; w[75][58] = 5'b00000; w[75][59] = 5'b01111; w[75][60] = 5'b01111; w[75][61] = 5'b01111; w[75][62] = 5'b00000; w[75][63] = 5'b10000; w[75][64] = 5'b01111; w[75][65] = 5'b01111; w[75][66] = 5'b01111; w[75][67] = 5'b00000; w[75][68] = 5'b01111; w[75][69] = 5'b01111; w[75][70] = 5'b01111; w[75][71] = 5'b01111; w[75][72] = 5'b00000; w[75][73] = 5'b01111; w[75][74] = 5'b01111; w[75][75] = 5'b00000; w[75][76] = 5'b00000; w[75][77] = 5'b10000; w[75][78] = 5'b01111; w[75][79] = 5'b01111; w[75][80] = 5'b01111; w[75][81] = 5'b00000; w[75][82] = 5'b01111; w[75][83] = 5'b01111; w[75][84] = 5'b01111; w[75][85] = 5'b01111; w[75][86] = 5'b00000; w[75][87] = 5'b01111; w[75][88] = 5'b01111; w[75][89] = 5'b01111; w[75][90] = 5'b00000; w[75][91] = 5'b00000; w[75][92] = 5'b01111; w[75][93] = 5'b01111; w[75][94] = 5'b01111; w[75][95] = 5'b01111; w[75][96] = 5'b01111; w[75][97] = 5'b01111; w[75][98] = 5'b01111; w[75][99] = 5'b01111; w[75][100] = 5'b00000; w[75][101] = 5'b01111; w[75][102] = 5'b01111; w[75][103] = 5'b01111; w[75][104] = 5'b00000; w[75][105] = 5'b00000; w[75][106] = 5'b00000; w[75][107] = 5'b01111; w[75][108] = 5'b01111; w[75][109] = 5'b00000; w[75][110] = 5'b01111; w[75][111] = 5'b01111; w[75][112] = 5'b01111; w[75][113] = 5'b01111; w[75][114] = 5'b00000; w[75][115] = 5'b01111; w[75][116] = 5'b01111; w[75][117] = 5'b01111; w[75][118] = 5'b00000; w[75][119] = 5'b00000; w[75][120] = 5'b01111; w[75][121] = 5'b01111; w[75][122] = 5'b01111; w[75][123] = 5'b00000; w[75][124] = 5'b01111; w[75][125] = 5'b01111; w[75][126] = 5'b01111; w[75][127] = 5'b01111; w[75][128] = 5'b00000; w[75][129] = 5'b01111; w[75][130] = 5'b01111; w[75][131] = 5'b01111; w[75][132] = 5'b10000; w[75][133] = 5'b00000; w[75][134] = 5'b01111; w[75][135] = 5'b01111; w[75][136] = 5'b01111; w[75][137] = 5'b00000; w[75][138] = 5'b01111; w[75][139] = 5'b01111; w[75][140] = 5'b01111; w[75][141] = 5'b01111; w[75][142] = 5'b00000; w[75][143] = 5'b01111; w[75][144] = 5'b01111; w[75][145] = 5'b01111; w[75][146] = 5'b10000; w[75][147] = 5'b00000; w[75][148] = 5'b01111; w[75][149] = 5'b01111; w[75][150] = 5'b01111; w[75][151] = 5'b00000; w[75][152] = 5'b01111; w[75][153] = 5'b01111; w[75][154] = 5'b01111; w[75][155] = 5'b01111; w[75][156] = 5'b01111; w[75][157] = 5'b01111; w[75][158] = 5'b01111; w[75][159] = 5'b10000; w[75][160] = 5'b10000; w[75][161] = 5'b10000; w[75][162] = 5'b00000; w[75][163] = 5'b01111; w[75][164] = 5'b01111; w[75][165] = 5'b01111; w[75][166] = 5'b01111; w[75][167] = 5'b01111; w[75][168] = 5'b01111; w[75][169] = 5'b01111; w[75][170] = 5'b01111; w[75][171] = 5'b01111; w[75][172] = 5'b01111; w[75][173] = 5'b10000; w[75][174] = 5'b10000; w[75][175] = 5'b10000; w[75][176] = 5'b00000; w[75][177] = 5'b01111; w[75][178] = 5'b01111; w[75][179] = 5'b01111; w[75][180] = 5'b01111; w[75][181] = 5'b01111; w[75][182] = 5'b01111; w[75][183] = 5'b01111; w[75][184] = 5'b01111; w[75][185] = 5'b01111; w[75][186] = 5'b01111; w[75][187] = 5'b01111; w[75][188] = 5'b01111; w[75][189] = 5'b01111; w[75][190] = 5'b01111; w[75][191] = 5'b01111; w[75][192] = 5'b01111; w[75][193] = 5'b01111; w[75][194] = 5'b01111; w[75][195] = 5'b01111; w[75][196] = 5'b01111; w[75][197] = 5'b01111; w[75][198] = 5'b01111; w[75][199] = 5'b01111; w[75][200] = 5'b01111; w[75][201] = 5'b01111; w[75][202] = 5'b01111; w[75][203] = 5'b01111; w[75][204] = 5'b01111; w[75][205] = 5'b01111; w[75][206] = 5'b01111; w[75][207] = 5'b01111; w[75][208] = 5'b01111; w[75][209] = 5'b01111; 
w[76][0] = 5'b10000; w[76][1] = 5'b10000; w[76][2] = 5'b10000; w[76][3] = 5'b10000; w[76][4] = 5'b10000; w[76][5] = 5'b10000; w[76][6] = 5'b10000; w[76][7] = 5'b10000; w[76][8] = 5'b10000; w[76][9] = 5'b10000; w[76][10] = 5'b10000; w[76][11] = 5'b10000; w[76][12] = 5'b10000; w[76][13] = 5'b10000; w[76][14] = 5'b10000; w[76][15] = 5'b10000; w[76][16] = 5'b10000; w[76][17] = 5'b10000; w[76][18] = 5'b10000; w[76][19] = 5'b10000; w[76][20] = 5'b10000; w[76][21] = 5'b10000; w[76][22] = 5'b10000; w[76][23] = 5'b10000; w[76][24] = 5'b10000; w[76][25] = 5'b10000; w[76][26] = 5'b10000; w[76][27] = 5'b10000; w[76][28] = 5'b10000; w[76][29] = 5'b10000; w[76][30] = 5'b00000; w[76][31] = 5'b01111; w[76][32] = 5'b00000; w[76][33] = 5'b01111; w[76][34] = 5'b00000; w[76][35] = 5'b00000; w[76][36] = 5'b00000; w[76][37] = 5'b00000; w[76][38] = 5'b01111; w[76][39] = 5'b00000; w[76][40] = 5'b10000; w[76][41] = 5'b10000; w[76][42] = 5'b10000; w[76][43] = 5'b10000; w[76][44] = 5'b00000; w[76][45] = 5'b00000; w[76][46] = 5'b00000; w[76][47] = 5'b01111; w[76][48] = 5'b00000; w[76][49] = 5'b00000; w[76][50] = 5'b00000; w[76][51] = 5'b00000; w[76][52] = 5'b00000; w[76][53] = 5'b00000; w[76][54] = 5'b10000; w[76][55] = 5'b10000; w[76][56] = 5'b10000; w[76][57] = 5'b10000; w[76][58] = 5'b10000; w[76][59] = 5'b10000; w[76][60] = 5'b10000; w[76][61] = 5'b00000; w[76][62] = 5'b01111; w[76][63] = 5'b01111; w[76][64] = 5'b10000; w[76][65] = 5'b10000; w[76][66] = 5'b10000; w[76][67] = 5'b10000; w[76][68] = 5'b10000; w[76][69] = 5'b10000; w[76][70] = 5'b10000; w[76][71] = 5'b10000; w[76][72] = 5'b10000; w[76][73] = 5'b10000; w[76][74] = 5'b00000; w[76][75] = 5'b00000; w[76][76] = 5'b00000; w[76][77] = 5'b01111; w[76][78] = 5'b10000; w[76][79] = 5'b00000; w[76][80] = 5'b10000; w[76][81] = 5'b10000; w[76][82] = 5'b10000; w[76][83] = 5'b10000; w[76][84] = 5'b10000; w[76][85] = 5'b10000; w[76][86] = 5'b10000; w[76][87] = 5'b10000; w[76][88] = 5'b00000; w[76][89] = 5'b00000; w[76][90] = 5'b01111; w[76][91] = 5'b01111; w[76][92] = 5'b10000; w[76][93] = 5'b00000; w[76][94] = 5'b00000; w[76][95] = 5'b10000; w[76][96] = 5'b10000; w[76][97] = 5'b10000; w[76][98] = 5'b10000; w[76][99] = 5'b10000; w[76][100] = 5'b10000; w[76][101] = 5'b10000; w[76][102] = 5'b00000; w[76][103] = 5'b10000; w[76][104] = 5'b01111; w[76][105] = 5'b01111; w[76][106] = 5'b10000; w[76][107] = 5'b10000; w[76][108] = 5'b10000; w[76][109] = 5'b10000; w[76][110] = 5'b10000; w[76][111] = 5'b10000; w[76][112] = 5'b10000; w[76][113] = 5'b10000; w[76][114] = 5'b10000; w[76][115] = 5'b10000; w[76][116] = 5'b00000; w[76][117] = 5'b10000; w[76][118] = 5'b01111; w[76][119] = 5'b01111; w[76][120] = 5'b10000; w[76][121] = 5'b10000; w[76][122] = 5'b10000; w[76][123] = 5'b10000; w[76][124] = 5'b10000; w[76][125] = 5'b10000; w[76][126] = 5'b10000; w[76][127] = 5'b10000; w[76][128] = 5'b10000; w[76][129] = 5'b10000; w[76][130] = 5'b00000; w[76][131] = 5'b10000; w[76][132] = 5'b01111; w[76][133] = 5'b01111; w[76][134] = 5'b00000; w[76][135] = 5'b00000; w[76][136] = 5'b10000; w[76][137] = 5'b10000; w[76][138] = 5'b10000; w[76][139] = 5'b10000; w[76][140] = 5'b10000; w[76][141] = 5'b10000; w[76][142] = 5'b10000; w[76][143] = 5'b10000; w[76][144] = 5'b10000; w[76][145] = 5'b10000; w[76][146] = 5'b01111; w[76][147] = 5'b01111; w[76][148] = 5'b00000; w[76][149] = 5'b10000; w[76][150] = 5'b10000; w[76][151] = 5'b10000; w[76][152] = 5'b10000; w[76][153] = 5'b10000; w[76][154] = 5'b10000; w[76][155] = 5'b10000; w[76][156] = 5'b10000; w[76][157] = 5'b10000; w[76][158] = 5'b10000; w[76][159] = 5'b10000; w[76][160] = 5'b00000; w[76][161] = 5'b00000; w[76][162] = 5'b00000; w[76][163] = 5'b10000; w[76][164] = 5'b10000; w[76][165] = 5'b10000; w[76][166] = 5'b10000; w[76][167] = 5'b10000; w[76][168] = 5'b10000; w[76][169] = 5'b10000; w[76][170] = 5'b10000; w[76][171] = 5'b00000; w[76][172] = 5'b10000; w[76][173] = 5'b10000; w[76][174] = 5'b00000; w[76][175] = 5'b00000; w[76][176] = 5'b00000; w[76][177] = 5'b10000; w[76][178] = 5'b00000; w[76][179] = 5'b10000; w[76][180] = 5'b10000; w[76][181] = 5'b10000; w[76][182] = 5'b10000; w[76][183] = 5'b10000; w[76][184] = 5'b10000; w[76][185] = 5'b10000; w[76][186] = 5'b10000; w[76][187] = 5'b10000; w[76][188] = 5'b10000; w[76][189] = 5'b10000; w[76][190] = 5'b10000; w[76][191] = 5'b10000; w[76][192] = 5'b10000; w[76][193] = 5'b10000; w[76][194] = 5'b10000; w[76][195] = 5'b10000; w[76][196] = 5'b10000; w[76][197] = 5'b10000; w[76][198] = 5'b10000; w[76][199] = 5'b10000; w[76][200] = 5'b10000; w[76][201] = 5'b10000; w[76][202] = 5'b10000; w[76][203] = 5'b10000; w[76][204] = 5'b10000; w[76][205] = 5'b10000; w[76][206] = 5'b10000; w[76][207] = 5'b10000; w[76][208] = 5'b10000; w[76][209] = 5'b10000; 
w[77][0] = 5'b00000; w[77][1] = 5'b00000; w[77][2] = 5'b00000; w[77][3] = 5'b00000; w[77][4] = 5'b00000; w[77][5] = 5'b00000; w[77][6] = 5'b00000; w[77][7] = 5'b00000; w[77][8] = 5'b00000; w[77][9] = 5'b00000; w[77][10] = 5'b00000; w[77][11] = 5'b00000; w[77][12] = 5'b00000; w[77][13] = 5'b00000; w[77][14] = 5'b00000; w[77][15] = 5'b00000; w[77][16] = 5'b00000; w[77][17] = 5'b00000; w[77][18] = 5'b00000; w[77][19] = 5'b00000; w[77][20] = 5'b00000; w[77][21] = 5'b00000; w[77][22] = 5'b00000; w[77][23] = 5'b00000; w[77][24] = 5'b00000; w[77][25] = 5'b00000; w[77][26] = 5'b00000; w[77][27] = 5'b00000; w[77][28] = 5'b00000; w[77][29] = 5'b00000; w[77][30] = 5'b01111; w[77][31] = 5'b00000; w[77][32] = 5'b10000; w[77][33] = 5'b00000; w[77][34] = 5'b01111; w[77][35] = 5'b01111; w[77][36] = 5'b01111; w[77][37] = 5'b10000; w[77][38] = 5'b00000; w[77][39] = 5'b01111; w[77][40] = 5'b00000; w[77][41] = 5'b00000; w[77][42] = 5'b00000; w[77][43] = 5'b00000; w[77][44] = 5'b01111; w[77][45] = 5'b10000; w[77][46] = 5'b10000; w[77][47] = 5'b00000; w[77][48] = 5'b01111; w[77][49] = 5'b01111; w[77][50] = 5'b01111; w[77][51] = 5'b10000; w[77][52] = 5'b10000; w[77][53] = 5'b01111; w[77][54] = 5'b00000; w[77][55] = 5'b00000; w[77][56] = 5'b00000; w[77][57] = 5'b00000; w[77][58] = 5'b10000; w[77][59] = 5'b10000; w[77][60] = 5'b10000; w[77][61] = 5'b10000; w[77][62] = 5'b01111; w[77][63] = 5'b01111; w[77][64] = 5'b00000; w[77][65] = 5'b10000; w[77][66] = 5'b10000; w[77][67] = 5'b10000; w[77][68] = 5'b00000; w[77][69] = 5'b00000; w[77][70] = 5'b00000; w[77][71] = 5'b00000; w[77][72] = 5'b10000; w[77][73] = 5'b10000; w[77][74] = 5'b10000; w[77][75] = 5'b10000; w[77][76] = 5'b01111; w[77][77] = 5'b00000; w[77][78] = 5'b00000; w[77][79] = 5'b10000; w[77][80] = 5'b10000; w[77][81] = 5'b10000; w[77][82] = 5'b00000; w[77][83] = 5'b00000; w[77][84] = 5'b00000; w[77][85] = 5'b00000; w[77][86] = 5'b10000; w[77][87] = 5'b10000; w[77][88] = 5'b10000; w[77][89] = 5'b10000; w[77][90] = 5'b01111; w[77][91] = 5'b01111; w[77][92] = 5'b00000; w[77][93] = 5'b10000; w[77][94] = 5'b10000; w[77][95] = 5'b00000; w[77][96] = 5'b00000; w[77][97] = 5'b00000; w[77][98] = 5'b00000; w[77][99] = 5'b00000; w[77][100] = 5'b10000; w[77][101] = 5'b10000; w[77][102] = 5'b10000; w[77][103] = 5'b00000; w[77][104] = 5'b01111; w[77][105] = 5'b01111; w[77][106] = 5'b10000; w[77][107] = 5'b10000; w[77][108] = 5'b10000; w[77][109] = 5'b10000; w[77][110] = 5'b00000; w[77][111] = 5'b00000; w[77][112] = 5'b00000; w[77][113] = 5'b00000; w[77][114] = 5'b10000; w[77][115] = 5'b10000; w[77][116] = 5'b10000; w[77][117] = 5'b00000; w[77][118] = 5'b01111; w[77][119] = 5'b01111; w[77][120] = 5'b10000; w[77][121] = 5'b10000; w[77][122] = 5'b10000; w[77][123] = 5'b10000; w[77][124] = 5'b00000; w[77][125] = 5'b00000; w[77][126] = 5'b00000; w[77][127] = 5'b00000; w[77][128] = 5'b10000; w[77][129] = 5'b10000; w[77][130] = 5'b10000; w[77][131] = 5'b00000; w[77][132] = 5'b01111; w[77][133] = 5'b01111; w[77][134] = 5'b10000; w[77][135] = 5'b10000; w[77][136] = 5'b10000; w[77][137] = 5'b10000; w[77][138] = 5'b00000; w[77][139] = 5'b00000; w[77][140] = 5'b00000; w[77][141] = 5'b00000; w[77][142] = 5'b10000; w[77][143] = 5'b10000; w[77][144] = 5'b10000; w[77][145] = 5'b00000; w[77][146] = 5'b01111; w[77][147] = 5'b01111; w[77][148] = 5'b10000; w[77][149] = 5'b10000; w[77][150] = 5'b10000; w[77][151] = 5'b10000; w[77][152] = 5'b00000; w[77][153] = 5'b00000; w[77][154] = 5'b00000; w[77][155] = 5'b00000; w[77][156] = 5'b00000; w[77][157] = 5'b10000; w[77][158] = 5'b10000; w[77][159] = 5'b00000; w[77][160] = 5'b01111; w[77][161] = 5'b01111; w[77][162] = 5'b10000; w[77][163] = 5'b10000; w[77][164] = 5'b10000; w[77][165] = 5'b00000; w[77][166] = 5'b00000; w[77][167] = 5'b00000; w[77][168] = 5'b00000; w[77][169] = 5'b00000; w[77][170] = 5'b00000; w[77][171] = 5'b10000; w[77][172] = 5'b10000; w[77][173] = 5'b00000; w[77][174] = 5'b01111; w[77][175] = 5'b01111; w[77][176] = 5'b10000; w[77][177] = 5'b10000; w[77][178] = 5'b10000; w[77][179] = 5'b00000; w[77][180] = 5'b00000; w[77][181] = 5'b00000; w[77][182] = 5'b00000; w[77][183] = 5'b00000; w[77][184] = 5'b00000; w[77][185] = 5'b00000; w[77][186] = 5'b00000; w[77][187] = 5'b00000; w[77][188] = 5'b00000; w[77][189] = 5'b00000; w[77][190] = 5'b00000; w[77][191] = 5'b00000; w[77][192] = 5'b00000; w[77][193] = 5'b00000; w[77][194] = 5'b00000; w[77][195] = 5'b00000; w[77][196] = 5'b00000; w[77][197] = 5'b00000; w[77][198] = 5'b00000; w[77][199] = 5'b00000; w[77][200] = 5'b00000; w[77][201] = 5'b00000; w[77][202] = 5'b00000; w[77][203] = 5'b00000; w[77][204] = 5'b00000; w[77][205] = 5'b00000; w[77][206] = 5'b00000; w[77][207] = 5'b00000; w[77][208] = 5'b00000; w[77][209] = 5'b00000; 
w[78][0] = 5'b01111; w[78][1] = 5'b01111; w[78][2] = 5'b01111; w[78][3] = 5'b01111; w[78][4] = 5'b01111; w[78][5] = 5'b01111; w[78][6] = 5'b01111; w[78][7] = 5'b01111; w[78][8] = 5'b01111; w[78][9] = 5'b01111; w[78][10] = 5'b01111; w[78][11] = 5'b01111; w[78][12] = 5'b01111; w[78][13] = 5'b01111; w[78][14] = 5'b01111; w[78][15] = 5'b01111; w[78][16] = 5'b01111; w[78][17] = 5'b01111; w[78][18] = 5'b01111; w[78][19] = 5'b01111; w[78][20] = 5'b01111; w[78][21] = 5'b01111; w[78][22] = 5'b01111; w[78][23] = 5'b01111; w[78][24] = 5'b01111; w[78][25] = 5'b01111; w[78][26] = 5'b01111; w[78][27] = 5'b01111; w[78][28] = 5'b01111; w[78][29] = 5'b01111; w[78][30] = 5'b01111; w[78][31] = 5'b00000; w[78][32] = 5'b10000; w[78][33] = 5'b10000; w[78][34] = 5'b10000; w[78][35] = 5'b10000; w[78][36] = 5'b10000; w[78][37] = 5'b10000; w[78][38] = 5'b00000; w[78][39] = 5'b01111; w[78][40] = 5'b01111; w[78][41] = 5'b01111; w[78][42] = 5'b01111; w[78][43] = 5'b01111; w[78][44] = 5'b01111; w[78][45] = 5'b10000; w[78][46] = 5'b10000; w[78][47] = 5'b10000; w[78][48] = 5'b10000; w[78][49] = 5'b10000; w[78][50] = 5'b10000; w[78][51] = 5'b10000; w[78][52] = 5'b10000; w[78][53] = 5'b01111; w[78][54] = 5'b01111; w[78][55] = 5'b01111; w[78][56] = 5'b01111; w[78][57] = 5'b01111; w[78][58] = 5'b01111; w[78][59] = 5'b00000; w[78][60] = 5'b00000; w[78][61] = 5'b01111; w[78][62] = 5'b10000; w[78][63] = 5'b00000; w[78][64] = 5'b01111; w[78][65] = 5'b00000; w[78][66] = 5'b00000; w[78][67] = 5'b01111; w[78][68] = 5'b01111; w[78][69] = 5'b01111; w[78][70] = 5'b01111; w[78][71] = 5'b01111; w[78][72] = 5'b01111; w[78][73] = 5'b00000; w[78][74] = 5'b01111; w[78][75] = 5'b01111; w[78][76] = 5'b10000; w[78][77] = 5'b00000; w[78][78] = 5'b00000; w[78][79] = 5'b01111; w[78][80] = 5'b00000; w[78][81] = 5'b01111; w[78][82] = 5'b01111; w[78][83] = 5'b01111; w[78][84] = 5'b01111; w[78][85] = 5'b01111; w[78][86] = 5'b01111; w[78][87] = 5'b00000; w[78][88] = 5'b01111; w[78][89] = 5'b01111; w[78][90] = 5'b10000; w[78][91] = 5'b10000; w[78][92] = 5'b01111; w[78][93] = 5'b01111; w[78][94] = 5'b01111; w[78][95] = 5'b01111; w[78][96] = 5'b01111; w[78][97] = 5'b01111; w[78][98] = 5'b01111; w[78][99] = 5'b01111; w[78][100] = 5'b01111; w[78][101] = 5'b00000; w[78][102] = 5'b01111; w[78][103] = 5'b01111; w[78][104] = 5'b10000; w[78][105] = 5'b10000; w[78][106] = 5'b01111; w[78][107] = 5'b00000; w[78][108] = 5'b00000; w[78][109] = 5'b01111; w[78][110] = 5'b01111; w[78][111] = 5'b01111; w[78][112] = 5'b01111; w[78][113] = 5'b01111; w[78][114] = 5'b01111; w[78][115] = 5'b00000; w[78][116] = 5'b01111; w[78][117] = 5'b01111; w[78][118] = 5'b10000; w[78][119] = 5'b10000; w[78][120] = 5'b00000; w[78][121] = 5'b00000; w[78][122] = 5'b00000; w[78][123] = 5'b01111; w[78][124] = 5'b01111; w[78][125] = 5'b01111; w[78][126] = 5'b01111; w[78][127] = 5'b01111; w[78][128] = 5'b01111; w[78][129] = 5'b00000; w[78][130] = 5'b01111; w[78][131] = 5'b01111; w[78][132] = 5'b00000; w[78][133] = 5'b10000; w[78][134] = 5'b01111; w[78][135] = 5'b01111; w[78][136] = 5'b00000; w[78][137] = 5'b01111; w[78][138] = 5'b01111; w[78][139] = 5'b01111; w[78][140] = 5'b01111; w[78][141] = 5'b01111; w[78][142] = 5'b01111; w[78][143] = 5'b00000; w[78][144] = 5'b00000; w[78][145] = 5'b01111; w[78][146] = 5'b00000; w[78][147] = 5'b10000; w[78][148] = 5'b01111; w[78][149] = 5'b00000; w[78][150] = 5'b00000; w[78][151] = 5'b01111; w[78][152] = 5'b01111; w[78][153] = 5'b01111; w[78][154] = 5'b01111; w[78][155] = 5'b01111; w[78][156] = 5'b01111; w[78][157] = 5'b00000; w[78][158] = 5'b00000; w[78][159] = 5'b00000; w[78][160] = 5'b10000; w[78][161] = 5'b10000; w[78][162] = 5'b10000; w[78][163] = 5'b00000; w[78][164] = 5'b00000; w[78][165] = 5'b01111; w[78][166] = 5'b01111; w[78][167] = 5'b01111; w[78][168] = 5'b01111; w[78][169] = 5'b01111; w[78][170] = 5'b01111; w[78][171] = 5'b01111; w[78][172] = 5'b00000; w[78][173] = 5'b00000; w[78][174] = 5'b10000; w[78][175] = 5'b10000; w[78][176] = 5'b10000; w[78][177] = 5'b00000; w[78][178] = 5'b01111; w[78][179] = 5'b01111; w[78][180] = 5'b01111; w[78][181] = 5'b01111; w[78][182] = 5'b01111; w[78][183] = 5'b01111; w[78][184] = 5'b01111; w[78][185] = 5'b01111; w[78][186] = 5'b01111; w[78][187] = 5'b01111; w[78][188] = 5'b01111; w[78][189] = 5'b01111; w[78][190] = 5'b01111; w[78][191] = 5'b01111; w[78][192] = 5'b01111; w[78][193] = 5'b01111; w[78][194] = 5'b01111; w[78][195] = 5'b01111; w[78][196] = 5'b01111; w[78][197] = 5'b01111; w[78][198] = 5'b01111; w[78][199] = 5'b01111; w[78][200] = 5'b01111; w[78][201] = 5'b01111; w[78][202] = 5'b01111; w[78][203] = 5'b01111; w[78][204] = 5'b01111; w[78][205] = 5'b01111; w[78][206] = 5'b01111; w[78][207] = 5'b01111; w[78][208] = 5'b01111; w[78][209] = 5'b01111; 
w[79][0] = 5'b01111; w[79][1] = 5'b01111; w[79][2] = 5'b01111; w[79][3] = 5'b01111; w[79][4] = 5'b01111; w[79][5] = 5'b01111; w[79][6] = 5'b01111; w[79][7] = 5'b01111; w[79][8] = 5'b01111; w[79][9] = 5'b01111; w[79][10] = 5'b01111; w[79][11] = 5'b01111; w[79][12] = 5'b01111; w[79][13] = 5'b01111; w[79][14] = 5'b01111; w[79][15] = 5'b01111; w[79][16] = 5'b01111; w[79][17] = 5'b01111; w[79][18] = 5'b01111; w[79][19] = 5'b01111; w[79][20] = 5'b01111; w[79][21] = 5'b01111; w[79][22] = 5'b01111; w[79][23] = 5'b01111; w[79][24] = 5'b01111; w[79][25] = 5'b01111; w[79][26] = 5'b01111; w[79][27] = 5'b01111; w[79][28] = 5'b01111; w[79][29] = 5'b01111; w[79][30] = 5'b00000; w[79][31] = 5'b01111; w[79][32] = 5'b00000; w[79][33] = 5'b10000; w[79][34] = 5'b10000; w[79][35] = 5'b10000; w[79][36] = 5'b10000; w[79][37] = 5'b00000; w[79][38] = 5'b01111; w[79][39] = 5'b00000; w[79][40] = 5'b01111; w[79][41] = 5'b01111; w[79][42] = 5'b01111; w[79][43] = 5'b01111; w[79][44] = 5'b00000; w[79][45] = 5'b00000; w[79][46] = 5'b00000; w[79][47] = 5'b10000; w[79][48] = 5'b10000; w[79][49] = 5'b10000; w[79][50] = 5'b10000; w[79][51] = 5'b00000; w[79][52] = 5'b00000; w[79][53] = 5'b00000; w[79][54] = 5'b01111; w[79][55] = 5'b01111; w[79][56] = 5'b01111; w[79][57] = 5'b01111; w[79][58] = 5'b00000; w[79][59] = 5'b01111; w[79][60] = 5'b01111; w[79][61] = 5'b01111; w[79][62] = 5'b00000; w[79][63] = 5'b10000; w[79][64] = 5'b01111; w[79][65] = 5'b01111; w[79][66] = 5'b01111; w[79][67] = 5'b00000; w[79][68] = 5'b01111; w[79][69] = 5'b01111; w[79][70] = 5'b01111; w[79][71] = 5'b01111; w[79][72] = 5'b00000; w[79][73] = 5'b01111; w[79][74] = 5'b01111; w[79][75] = 5'b01111; w[79][76] = 5'b00000; w[79][77] = 5'b10000; w[79][78] = 5'b01111; w[79][79] = 5'b00000; w[79][80] = 5'b01111; w[79][81] = 5'b00000; w[79][82] = 5'b01111; w[79][83] = 5'b01111; w[79][84] = 5'b01111; w[79][85] = 5'b01111; w[79][86] = 5'b00000; w[79][87] = 5'b01111; w[79][88] = 5'b01111; w[79][89] = 5'b01111; w[79][90] = 5'b00000; w[79][91] = 5'b00000; w[79][92] = 5'b01111; w[79][93] = 5'b01111; w[79][94] = 5'b01111; w[79][95] = 5'b01111; w[79][96] = 5'b01111; w[79][97] = 5'b01111; w[79][98] = 5'b01111; w[79][99] = 5'b01111; w[79][100] = 5'b00000; w[79][101] = 5'b01111; w[79][102] = 5'b01111; w[79][103] = 5'b01111; w[79][104] = 5'b00000; w[79][105] = 5'b00000; w[79][106] = 5'b00000; w[79][107] = 5'b01111; w[79][108] = 5'b01111; w[79][109] = 5'b00000; w[79][110] = 5'b01111; w[79][111] = 5'b01111; w[79][112] = 5'b01111; w[79][113] = 5'b01111; w[79][114] = 5'b00000; w[79][115] = 5'b01111; w[79][116] = 5'b01111; w[79][117] = 5'b01111; w[79][118] = 5'b00000; w[79][119] = 5'b00000; w[79][120] = 5'b01111; w[79][121] = 5'b01111; w[79][122] = 5'b01111; w[79][123] = 5'b00000; w[79][124] = 5'b01111; w[79][125] = 5'b01111; w[79][126] = 5'b01111; w[79][127] = 5'b01111; w[79][128] = 5'b00000; w[79][129] = 5'b01111; w[79][130] = 5'b01111; w[79][131] = 5'b01111; w[79][132] = 5'b10000; w[79][133] = 5'b00000; w[79][134] = 5'b01111; w[79][135] = 5'b01111; w[79][136] = 5'b01111; w[79][137] = 5'b00000; w[79][138] = 5'b01111; w[79][139] = 5'b01111; w[79][140] = 5'b01111; w[79][141] = 5'b01111; w[79][142] = 5'b00000; w[79][143] = 5'b01111; w[79][144] = 5'b01111; w[79][145] = 5'b01111; w[79][146] = 5'b10000; w[79][147] = 5'b00000; w[79][148] = 5'b01111; w[79][149] = 5'b01111; w[79][150] = 5'b01111; w[79][151] = 5'b00000; w[79][152] = 5'b01111; w[79][153] = 5'b01111; w[79][154] = 5'b01111; w[79][155] = 5'b01111; w[79][156] = 5'b01111; w[79][157] = 5'b01111; w[79][158] = 5'b01111; w[79][159] = 5'b10000; w[79][160] = 5'b10000; w[79][161] = 5'b10000; w[79][162] = 5'b00000; w[79][163] = 5'b01111; w[79][164] = 5'b01111; w[79][165] = 5'b01111; w[79][166] = 5'b01111; w[79][167] = 5'b01111; w[79][168] = 5'b01111; w[79][169] = 5'b01111; w[79][170] = 5'b01111; w[79][171] = 5'b01111; w[79][172] = 5'b01111; w[79][173] = 5'b10000; w[79][174] = 5'b10000; w[79][175] = 5'b10000; w[79][176] = 5'b00000; w[79][177] = 5'b01111; w[79][178] = 5'b01111; w[79][179] = 5'b01111; w[79][180] = 5'b01111; w[79][181] = 5'b01111; w[79][182] = 5'b01111; w[79][183] = 5'b01111; w[79][184] = 5'b01111; w[79][185] = 5'b01111; w[79][186] = 5'b01111; w[79][187] = 5'b01111; w[79][188] = 5'b01111; w[79][189] = 5'b01111; w[79][190] = 5'b01111; w[79][191] = 5'b01111; w[79][192] = 5'b01111; w[79][193] = 5'b01111; w[79][194] = 5'b01111; w[79][195] = 5'b01111; w[79][196] = 5'b01111; w[79][197] = 5'b01111; w[79][198] = 5'b01111; w[79][199] = 5'b01111; w[79][200] = 5'b01111; w[79][201] = 5'b01111; w[79][202] = 5'b01111; w[79][203] = 5'b01111; w[79][204] = 5'b01111; w[79][205] = 5'b01111; w[79][206] = 5'b01111; w[79][207] = 5'b01111; w[79][208] = 5'b01111; w[79][209] = 5'b01111; 
w[80][0] = 5'b00000; w[80][1] = 5'b00000; w[80][2] = 5'b00000; w[80][3] = 5'b00000; w[80][4] = 5'b00000; w[80][5] = 5'b00000; w[80][6] = 5'b00000; w[80][7] = 5'b00000; w[80][8] = 5'b00000; w[80][9] = 5'b00000; w[80][10] = 5'b00000; w[80][11] = 5'b00000; w[80][12] = 5'b00000; w[80][13] = 5'b00000; w[80][14] = 5'b00000; w[80][15] = 5'b00000; w[80][16] = 5'b00000; w[80][17] = 5'b00000; w[80][18] = 5'b00000; w[80][19] = 5'b00000; w[80][20] = 5'b00000; w[80][21] = 5'b00000; w[80][22] = 5'b00000; w[80][23] = 5'b00000; w[80][24] = 5'b00000; w[80][25] = 5'b00000; w[80][26] = 5'b00000; w[80][27] = 5'b00000; w[80][28] = 5'b00000; w[80][29] = 5'b00000; w[80][30] = 5'b10000; w[80][31] = 5'b00000; w[80][32] = 5'b01111; w[80][33] = 5'b00000; w[80][34] = 5'b10000; w[80][35] = 5'b10000; w[80][36] = 5'b10000; w[80][37] = 5'b01111; w[80][38] = 5'b00000; w[80][39] = 5'b10000; w[80][40] = 5'b00000; w[80][41] = 5'b00000; w[80][42] = 5'b00000; w[80][43] = 5'b00000; w[80][44] = 5'b10000; w[80][45] = 5'b01111; w[80][46] = 5'b01111; w[80][47] = 5'b00000; w[80][48] = 5'b10000; w[80][49] = 5'b10000; w[80][50] = 5'b10000; w[80][51] = 5'b01111; w[80][52] = 5'b01111; w[80][53] = 5'b10000; w[80][54] = 5'b00000; w[80][55] = 5'b00000; w[80][56] = 5'b00000; w[80][57] = 5'b00000; w[80][58] = 5'b01111; w[80][59] = 5'b01111; w[80][60] = 5'b01111; w[80][61] = 5'b01111; w[80][62] = 5'b10000; w[80][63] = 5'b10000; w[80][64] = 5'b00000; w[80][65] = 5'b01111; w[80][66] = 5'b01111; w[80][67] = 5'b01111; w[80][68] = 5'b00000; w[80][69] = 5'b00000; w[80][70] = 5'b00000; w[80][71] = 5'b00000; w[80][72] = 5'b01111; w[80][73] = 5'b01111; w[80][74] = 5'b01111; w[80][75] = 5'b01111; w[80][76] = 5'b10000; w[80][77] = 5'b10000; w[80][78] = 5'b00000; w[80][79] = 5'b01111; w[80][80] = 5'b00000; w[80][81] = 5'b01111; w[80][82] = 5'b00000; w[80][83] = 5'b00000; w[80][84] = 5'b00000; w[80][85] = 5'b00000; w[80][86] = 5'b01111; w[80][87] = 5'b01111; w[80][88] = 5'b01111; w[80][89] = 5'b01111; w[80][90] = 5'b10000; w[80][91] = 5'b10000; w[80][92] = 5'b00000; w[80][93] = 5'b01111; w[80][94] = 5'b01111; w[80][95] = 5'b00000; w[80][96] = 5'b00000; w[80][97] = 5'b00000; w[80][98] = 5'b00000; w[80][99] = 5'b00000; w[80][100] = 5'b01111; w[80][101] = 5'b01111; w[80][102] = 5'b01111; w[80][103] = 5'b00000; w[80][104] = 5'b10000; w[80][105] = 5'b10000; w[80][106] = 5'b01111; w[80][107] = 5'b01111; w[80][108] = 5'b01111; w[80][109] = 5'b01111; w[80][110] = 5'b00000; w[80][111] = 5'b00000; w[80][112] = 5'b00000; w[80][113] = 5'b00000; w[80][114] = 5'b01111; w[80][115] = 5'b01111; w[80][116] = 5'b01111; w[80][117] = 5'b00000; w[80][118] = 5'b10000; w[80][119] = 5'b10000; w[80][120] = 5'b01111; w[80][121] = 5'b01111; w[80][122] = 5'b01111; w[80][123] = 5'b01111; w[80][124] = 5'b00000; w[80][125] = 5'b00000; w[80][126] = 5'b00000; w[80][127] = 5'b00000; w[80][128] = 5'b01111; w[80][129] = 5'b01111; w[80][130] = 5'b01111; w[80][131] = 5'b00000; w[80][132] = 5'b10000; w[80][133] = 5'b10000; w[80][134] = 5'b01111; w[80][135] = 5'b01111; w[80][136] = 5'b01111; w[80][137] = 5'b01111; w[80][138] = 5'b00000; w[80][139] = 5'b00000; w[80][140] = 5'b00000; w[80][141] = 5'b00000; w[80][142] = 5'b01111; w[80][143] = 5'b01111; w[80][144] = 5'b01111; w[80][145] = 5'b00000; w[80][146] = 5'b10000; w[80][147] = 5'b10000; w[80][148] = 5'b01111; w[80][149] = 5'b01111; w[80][150] = 5'b01111; w[80][151] = 5'b01111; w[80][152] = 5'b00000; w[80][153] = 5'b00000; w[80][154] = 5'b00000; w[80][155] = 5'b00000; w[80][156] = 5'b00000; w[80][157] = 5'b01111; w[80][158] = 5'b01111; w[80][159] = 5'b00000; w[80][160] = 5'b10000; w[80][161] = 5'b10000; w[80][162] = 5'b01111; w[80][163] = 5'b01111; w[80][164] = 5'b01111; w[80][165] = 5'b00000; w[80][166] = 5'b00000; w[80][167] = 5'b00000; w[80][168] = 5'b00000; w[80][169] = 5'b00000; w[80][170] = 5'b00000; w[80][171] = 5'b01111; w[80][172] = 5'b01111; w[80][173] = 5'b00000; w[80][174] = 5'b10000; w[80][175] = 5'b10000; w[80][176] = 5'b01111; w[80][177] = 5'b01111; w[80][178] = 5'b01111; w[80][179] = 5'b00000; w[80][180] = 5'b00000; w[80][181] = 5'b00000; w[80][182] = 5'b00000; w[80][183] = 5'b00000; w[80][184] = 5'b00000; w[80][185] = 5'b00000; w[80][186] = 5'b00000; w[80][187] = 5'b00000; w[80][188] = 5'b00000; w[80][189] = 5'b00000; w[80][190] = 5'b00000; w[80][191] = 5'b00000; w[80][192] = 5'b00000; w[80][193] = 5'b00000; w[80][194] = 5'b00000; w[80][195] = 5'b00000; w[80][196] = 5'b00000; w[80][197] = 5'b00000; w[80][198] = 5'b00000; w[80][199] = 5'b00000; w[80][200] = 5'b00000; w[80][201] = 5'b00000; w[80][202] = 5'b00000; w[80][203] = 5'b00000; w[80][204] = 5'b00000; w[80][205] = 5'b00000; w[80][206] = 5'b00000; w[80][207] = 5'b00000; w[80][208] = 5'b00000; w[80][209] = 5'b00000; 
w[81][0] = 5'b01111; w[81][1] = 5'b01111; w[81][2] = 5'b01111; w[81][3] = 5'b01111; w[81][4] = 5'b01111; w[81][5] = 5'b01111; w[81][6] = 5'b01111; w[81][7] = 5'b01111; w[81][8] = 5'b01111; w[81][9] = 5'b01111; w[81][10] = 5'b01111; w[81][11] = 5'b01111; w[81][12] = 5'b01111; w[81][13] = 5'b01111; w[81][14] = 5'b01111; w[81][15] = 5'b01111; w[81][16] = 5'b01111; w[81][17] = 5'b01111; w[81][18] = 5'b01111; w[81][19] = 5'b01111; w[81][20] = 5'b01111; w[81][21] = 5'b01111; w[81][22] = 5'b01111; w[81][23] = 5'b01111; w[81][24] = 5'b01111; w[81][25] = 5'b01111; w[81][26] = 5'b01111; w[81][27] = 5'b01111; w[81][28] = 5'b01111; w[81][29] = 5'b01111; w[81][30] = 5'b00000; w[81][31] = 5'b10000; w[81][32] = 5'b00000; w[81][33] = 5'b10000; w[81][34] = 5'b00000; w[81][35] = 5'b00000; w[81][36] = 5'b00000; w[81][37] = 5'b00000; w[81][38] = 5'b10000; w[81][39] = 5'b00000; w[81][40] = 5'b01111; w[81][41] = 5'b01111; w[81][42] = 5'b01111; w[81][43] = 5'b01111; w[81][44] = 5'b00000; w[81][45] = 5'b00000; w[81][46] = 5'b00000; w[81][47] = 5'b10000; w[81][48] = 5'b00000; w[81][49] = 5'b00000; w[81][50] = 5'b00000; w[81][51] = 5'b00000; w[81][52] = 5'b00000; w[81][53] = 5'b00000; w[81][54] = 5'b01111; w[81][55] = 5'b01111; w[81][56] = 5'b01111; w[81][57] = 5'b01111; w[81][58] = 5'b01111; w[81][59] = 5'b01111; w[81][60] = 5'b01111; w[81][61] = 5'b00000; w[81][62] = 5'b10000; w[81][63] = 5'b10000; w[81][64] = 5'b01111; w[81][65] = 5'b01111; w[81][66] = 5'b01111; w[81][67] = 5'b01111; w[81][68] = 5'b01111; w[81][69] = 5'b01111; w[81][70] = 5'b01111; w[81][71] = 5'b01111; w[81][72] = 5'b01111; w[81][73] = 5'b01111; w[81][74] = 5'b00000; w[81][75] = 5'b00000; w[81][76] = 5'b10000; w[81][77] = 5'b10000; w[81][78] = 5'b01111; w[81][79] = 5'b00000; w[81][80] = 5'b01111; w[81][81] = 5'b00000; w[81][82] = 5'b01111; w[81][83] = 5'b01111; w[81][84] = 5'b01111; w[81][85] = 5'b01111; w[81][86] = 5'b01111; w[81][87] = 5'b01111; w[81][88] = 5'b00000; w[81][89] = 5'b00000; w[81][90] = 5'b10000; w[81][91] = 5'b10000; w[81][92] = 5'b01111; w[81][93] = 5'b00000; w[81][94] = 5'b00000; w[81][95] = 5'b01111; w[81][96] = 5'b01111; w[81][97] = 5'b01111; w[81][98] = 5'b01111; w[81][99] = 5'b01111; w[81][100] = 5'b01111; w[81][101] = 5'b01111; w[81][102] = 5'b00000; w[81][103] = 5'b01111; w[81][104] = 5'b10000; w[81][105] = 5'b10000; w[81][106] = 5'b01111; w[81][107] = 5'b01111; w[81][108] = 5'b01111; w[81][109] = 5'b01111; w[81][110] = 5'b01111; w[81][111] = 5'b01111; w[81][112] = 5'b01111; w[81][113] = 5'b01111; w[81][114] = 5'b01111; w[81][115] = 5'b01111; w[81][116] = 5'b00000; w[81][117] = 5'b01111; w[81][118] = 5'b10000; w[81][119] = 5'b10000; w[81][120] = 5'b01111; w[81][121] = 5'b01111; w[81][122] = 5'b01111; w[81][123] = 5'b01111; w[81][124] = 5'b01111; w[81][125] = 5'b01111; w[81][126] = 5'b01111; w[81][127] = 5'b01111; w[81][128] = 5'b01111; w[81][129] = 5'b01111; w[81][130] = 5'b00000; w[81][131] = 5'b01111; w[81][132] = 5'b10000; w[81][133] = 5'b10000; w[81][134] = 5'b00000; w[81][135] = 5'b00000; w[81][136] = 5'b01111; w[81][137] = 5'b01111; w[81][138] = 5'b01111; w[81][139] = 5'b01111; w[81][140] = 5'b01111; w[81][141] = 5'b01111; w[81][142] = 5'b01111; w[81][143] = 5'b01111; w[81][144] = 5'b01111; w[81][145] = 5'b01111; w[81][146] = 5'b10000; w[81][147] = 5'b10000; w[81][148] = 5'b00000; w[81][149] = 5'b01111; w[81][150] = 5'b01111; w[81][151] = 5'b01111; w[81][152] = 5'b01111; w[81][153] = 5'b01111; w[81][154] = 5'b01111; w[81][155] = 5'b01111; w[81][156] = 5'b01111; w[81][157] = 5'b01111; w[81][158] = 5'b01111; w[81][159] = 5'b01111; w[81][160] = 5'b00000; w[81][161] = 5'b00000; w[81][162] = 5'b00000; w[81][163] = 5'b01111; w[81][164] = 5'b01111; w[81][165] = 5'b01111; w[81][166] = 5'b01111; w[81][167] = 5'b01111; w[81][168] = 5'b01111; w[81][169] = 5'b01111; w[81][170] = 5'b01111; w[81][171] = 5'b00000; w[81][172] = 5'b01111; w[81][173] = 5'b01111; w[81][174] = 5'b00000; w[81][175] = 5'b00000; w[81][176] = 5'b00000; w[81][177] = 5'b01111; w[81][178] = 5'b00000; w[81][179] = 5'b01111; w[81][180] = 5'b01111; w[81][181] = 5'b01111; w[81][182] = 5'b01111; w[81][183] = 5'b01111; w[81][184] = 5'b01111; w[81][185] = 5'b01111; w[81][186] = 5'b01111; w[81][187] = 5'b01111; w[81][188] = 5'b01111; w[81][189] = 5'b01111; w[81][190] = 5'b01111; w[81][191] = 5'b01111; w[81][192] = 5'b01111; w[81][193] = 5'b01111; w[81][194] = 5'b01111; w[81][195] = 5'b01111; w[81][196] = 5'b01111; w[81][197] = 5'b01111; w[81][198] = 5'b01111; w[81][199] = 5'b01111; w[81][200] = 5'b01111; w[81][201] = 5'b01111; w[81][202] = 5'b01111; w[81][203] = 5'b01111; w[81][204] = 5'b01111; w[81][205] = 5'b01111; w[81][206] = 5'b01111; w[81][207] = 5'b01111; w[81][208] = 5'b01111; w[81][209] = 5'b01111; 
w[82][0] = 5'b01111; w[82][1] = 5'b01111; w[82][2] = 5'b01111; w[82][3] = 5'b01111; w[82][4] = 5'b01111; w[82][5] = 5'b01111; w[82][6] = 5'b01111; w[82][7] = 5'b01111; w[82][8] = 5'b01111; w[82][9] = 5'b01111; w[82][10] = 5'b01111; w[82][11] = 5'b01111; w[82][12] = 5'b01111; w[82][13] = 5'b01111; w[82][14] = 5'b01111; w[82][15] = 5'b01111; w[82][16] = 5'b01111; w[82][17] = 5'b01111; w[82][18] = 5'b01111; w[82][19] = 5'b01111; w[82][20] = 5'b01111; w[82][21] = 5'b01111; w[82][22] = 5'b01111; w[82][23] = 5'b01111; w[82][24] = 5'b01111; w[82][25] = 5'b01111; w[82][26] = 5'b01111; w[82][27] = 5'b01111; w[82][28] = 5'b01111; w[82][29] = 5'b01111; w[82][30] = 5'b01111; w[82][31] = 5'b00000; w[82][32] = 5'b10000; w[82][33] = 5'b10000; w[82][34] = 5'b10000; w[82][35] = 5'b10000; w[82][36] = 5'b10000; w[82][37] = 5'b10000; w[82][38] = 5'b00000; w[82][39] = 5'b01111; w[82][40] = 5'b01111; w[82][41] = 5'b01111; w[82][42] = 5'b01111; w[82][43] = 5'b01111; w[82][44] = 5'b01111; w[82][45] = 5'b10000; w[82][46] = 5'b10000; w[82][47] = 5'b10000; w[82][48] = 5'b10000; w[82][49] = 5'b10000; w[82][50] = 5'b10000; w[82][51] = 5'b10000; w[82][52] = 5'b10000; w[82][53] = 5'b01111; w[82][54] = 5'b01111; w[82][55] = 5'b01111; w[82][56] = 5'b01111; w[82][57] = 5'b01111; w[82][58] = 5'b01111; w[82][59] = 5'b00000; w[82][60] = 5'b00000; w[82][61] = 5'b01111; w[82][62] = 5'b10000; w[82][63] = 5'b00000; w[82][64] = 5'b01111; w[82][65] = 5'b00000; w[82][66] = 5'b00000; w[82][67] = 5'b01111; w[82][68] = 5'b01111; w[82][69] = 5'b01111; w[82][70] = 5'b01111; w[82][71] = 5'b01111; w[82][72] = 5'b01111; w[82][73] = 5'b00000; w[82][74] = 5'b01111; w[82][75] = 5'b01111; w[82][76] = 5'b10000; w[82][77] = 5'b00000; w[82][78] = 5'b01111; w[82][79] = 5'b01111; w[82][80] = 5'b00000; w[82][81] = 5'b01111; w[82][82] = 5'b00000; w[82][83] = 5'b01111; w[82][84] = 5'b01111; w[82][85] = 5'b01111; w[82][86] = 5'b01111; w[82][87] = 5'b00000; w[82][88] = 5'b01111; w[82][89] = 5'b01111; w[82][90] = 5'b10000; w[82][91] = 5'b10000; w[82][92] = 5'b01111; w[82][93] = 5'b01111; w[82][94] = 5'b01111; w[82][95] = 5'b01111; w[82][96] = 5'b01111; w[82][97] = 5'b01111; w[82][98] = 5'b01111; w[82][99] = 5'b01111; w[82][100] = 5'b01111; w[82][101] = 5'b00000; w[82][102] = 5'b01111; w[82][103] = 5'b01111; w[82][104] = 5'b10000; w[82][105] = 5'b10000; w[82][106] = 5'b01111; w[82][107] = 5'b00000; w[82][108] = 5'b00000; w[82][109] = 5'b01111; w[82][110] = 5'b01111; w[82][111] = 5'b01111; w[82][112] = 5'b01111; w[82][113] = 5'b01111; w[82][114] = 5'b01111; w[82][115] = 5'b00000; w[82][116] = 5'b01111; w[82][117] = 5'b01111; w[82][118] = 5'b10000; w[82][119] = 5'b10000; w[82][120] = 5'b00000; w[82][121] = 5'b00000; w[82][122] = 5'b00000; w[82][123] = 5'b01111; w[82][124] = 5'b01111; w[82][125] = 5'b01111; w[82][126] = 5'b01111; w[82][127] = 5'b01111; w[82][128] = 5'b01111; w[82][129] = 5'b00000; w[82][130] = 5'b01111; w[82][131] = 5'b01111; w[82][132] = 5'b00000; w[82][133] = 5'b10000; w[82][134] = 5'b01111; w[82][135] = 5'b01111; w[82][136] = 5'b00000; w[82][137] = 5'b01111; w[82][138] = 5'b01111; w[82][139] = 5'b01111; w[82][140] = 5'b01111; w[82][141] = 5'b01111; w[82][142] = 5'b01111; w[82][143] = 5'b00000; w[82][144] = 5'b00000; w[82][145] = 5'b01111; w[82][146] = 5'b00000; w[82][147] = 5'b10000; w[82][148] = 5'b01111; w[82][149] = 5'b00000; w[82][150] = 5'b00000; w[82][151] = 5'b01111; w[82][152] = 5'b01111; w[82][153] = 5'b01111; w[82][154] = 5'b01111; w[82][155] = 5'b01111; w[82][156] = 5'b01111; w[82][157] = 5'b00000; w[82][158] = 5'b00000; w[82][159] = 5'b00000; w[82][160] = 5'b10000; w[82][161] = 5'b10000; w[82][162] = 5'b10000; w[82][163] = 5'b00000; w[82][164] = 5'b00000; w[82][165] = 5'b01111; w[82][166] = 5'b01111; w[82][167] = 5'b01111; w[82][168] = 5'b01111; w[82][169] = 5'b01111; w[82][170] = 5'b01111; w[82][171] = 5'b01111; w[82][172] = 5'b00000; w[82][173] = 5'b00000; w[82][174] = 5'b10000; w[82][175] = 5'b10000; w[82][176] = 5'b10000; w[82][177] = 5'b00000; w[82][178] = 5'b01111; w[82][179] = 5'b01111; w[82][180] = 5'b01111; w[82][181] = 5'b01111; w[82][182] = 5'b01111; w[82][183] = 5'b01111; w[82][184] = 5'b01111; w[82][185] = 5'b01111; w[82][186] = 5'b01111; w[82][187] = 5'b01111; w[82][188] = 5'b01111; w[82][189] = 5'b01111; w[82][190] = 5'b01111; w[82][191] = 5'b01111; w[82][192] = 5'b01111; w[82][193] = 5'b01111; w[82][194] = 5'b01111; w[82][195] = 5'b01111; w[82][196] = 5'b01111; w[82][197] = 5'b01111; w[82][198] = 5'b01111; w[82][199] = 5'b01111; w[82][200] = 5'b01111; w[82][201] = 5'b01111; w[82][202] = 5'b01111; w[82][203] = 5'b01111; w[82][204] = 5'b01111; w[82][205] = 5'b01111; w[82][206] = 5'b01111; w[82][207] = 5'b01111; w[82][208] = 5'b01111; w[82][209] = 5'b01111; 
w[83][0] = 5'b01111; w[83][1] = 5'b01111; w[83][2] = 5'b01111; w[83][3] = 5'b01111; w[83][4] = 5'b01111; w[83][5] = 5'b01111; w[83][6] = 5'b01111; w[83][7] = 5'b01111; w[83][8] = 5'b01111; w[83][9] = 5'b01111; w[83][10] = 5'b01111; w[83][11] = 5'b01111; w[83][12] = 5'b01111; w[83][13] = 5'b01111; w[83][14] = 5'b01111; w[83][15] = 5'b01111; w[83][16] = 5'b01111; w[83][17] = 5'b01111; w[83][18] = 5'b01111; w[83][19] = 5'b01111; w[83][20] = 5'b01111; w[83][21] = 5'b01111; w[83][22] = 5'b01111; w[83][23] = 5'b01111; w[83][24] = 5'b01111; w[83][25] = 5'b01111; w[83][26] = 5'b01111; w[83][27] = 5'b01111; w[83][28] = 5'b01111; w[83][29] = 5'b01111; w[83][30] = 5'b01111; w[83][31] = 5'b00000; w[83][32] = 5'b10000; w[83][33] = 5'b10000; w[83][34] = 5'b10000; w[83][35] = 5'b10000; w[83][36] = 5'b10000; w[83][37] = 5'b10000; w[83][38] = 5'b00000; w[83][39] = 5'b01111; w[83][40] = 5'b01111; w[83][41] = 5'b01111; w[83][42] = 5'b01111; w[83][43] = 5'b01111; w[83][44] = 5'b01111; w[83][45] = 5'b10000; w[83][46] = 5'b10000; w[83][47] = 5'b10000; w[83][48] = 5'b10000; w[83][49] = 5'b10000; w[83][50] = 5'b10000; w[83][51] = 5'b10000; w[83][52] = 5'b10000; w[83][53] = 5'b01111; w[83][54] = 5'b01111; w[83][55] = 5'b01111; w[83][56] = 5'b01111; w[83][57] = 5'b01111; w[83][58] = 5'b01111; w[83][59] = 5'b00000; w[83][60] = 5'b00000; w[83][61] = 5'b01111; w[83][62] = 5'b10000; w[83][63] = 5'b00000; w[83][64] = 5'b01111; w[83][65] = 5'b00000; w[83][66] = 5'b00000; w[83][67] = 5'b01111; w[83][68] = 5'b01111; w[83][69] = 5'b01111; w[83][70] = 5'b01111; w[83][71] = 5'b01111; w[83][72] = 5'b01111; w[83][73] = 5'b00000; w[83][74] = 5'b01111; w[83][75] = 5'b01111; w[83][76] = 5'b10000; w[83][77] = 5'b00000; w[83][78] = 5'b01111; w[83][79] = 5'b01111; w[83][80] = 5'b00000; w[83][81] = 5'b01111; w[83][82] = 5'b01111; w[83][83] = 5'b00000; w[83][84] = 5'b01111; w[83][85] = 5'b01111; w[83][86] = 5'b01111; w[83][87] = 5'b00000; w[83][88] = 5'b01111; w[83][89] = 5'b01111; w[83][90] = 5'b10000; w[83][91] = 5'b10000; w[83][92] = 5'b01111; w[83][93] = 5'b01111; w[83][94] = 5'b01111; w[83][95] = 5'b01111; w[83][96] = 5'b01111; w[83][97] = 5'b01111; w[83][98] = 5'b01111; w[83][99] = 5'b01111; w[83][100] = 5'b01111; w[83][101] = 5'b00000; w[83][102] = 5'b01111; w[83][103] = 5'b01111; w[83][104] = 5'b10000; w[83][105] = 5'b10000; w[83][106] = 5'b01111; w[83][107] = 5'b00000; w[83][108] = 5'b00000; w[83][109] = 5'b01111; w[83][110] = 5'b01111; w[83][111] = 5'b01111; w[83][112] = 5'b01111; w[83][113] = 5'b01111; w[83][114] = 5'b01111; w[83][115] = 5'b00000; w[83][116] = 5'b01111; w[83][117] = 5'b01111; w[83][118] = 5'b10000; w[83][119] = 5'b10000; w[83][120] = 5'b00000; w[83][121] = 5'b00000; w[83][122] = 5'b00000; w[83][123] = 5'b01111; w[83][124] = 5'b01111; w[83][125] = 5'b01111; w[83][126] = 5'b01111; w[83][127] = 5'b01111; w[83][128] = 5'b01111; w[83][129] = 5'b00000; w[83][130] = 5'b01111; w[83][131] = 5'b01111; w[83][132] = 5'b00000; w[83][133] = 5'b10000; w[83][134] = 5'b01111; w[83][135] = 5'b01111; w[83][136] = 5'b00000; w[83][137] = 5'b01111; w[83][138] = 5'b01111; w[83][139] = 5'b01111; w[83][140] = 5'b01111; w[83][141] = 5'b01111; w[83][142] = 5'b01111; w[83][143] = 5'b00000; w[83][144] = 5'b00000; w[83][145] = 5'b01111; w[83][146] = 5'b00000; w[83][147] = 5'b10000; w[83][148] = 5'b01111; w[83][149] = 5'b00000; w[83][150] = 5'b00000; w[83][151] = 5'b01111; w[83][152] = 5'b01111; w[83][153] = 5'b01111; w[83][154] = 5'b01111; w[83][155] = 5'b01111; w[83][156] = 5'b01111; w[83][157] = 5'b00000; w[83][158] = 5'b00000; w[83][159] = 5'b00000; w[83][160] = 5'b10000; w[83][161] = 5'b10000; w[83][162] = 5'b10000; w[83][163] = 5'b00000; w[83][164] = 5'b00000; w[83][165] = 5'b01111; w[83][166] = 5'b01111; w[83][167] = 5'b01111; w[83][168] = 5'b01111; w[83][169] = 5'b01111; w[83][170] = 5'b01111; w[83][171] = 5'b01111; w[83][172] = 5'b00000; w[83][173] = 5'b00000; w[83][174] = 5'b10000; w[83][175] = 5'b10000; w[83][176] = 5'b10000; w[83][177] = 5'b00000; w[83][178] = 5'b01111; w[83][179] = 5'b01111; w[83][180] = 5'b01111; w[83][181] = 5'b01111; w[83][182] = 5'b01111; w[83][183] = 5'b01111; w[83][184] = 5'b01111; w[83][185] = 5'b01111; w[83][186] = 5'b01111; w[83][187] = 5'b01111; w[83][188] = 5'b01111; w[83][189] = 5'b01111; w[83][190] = 5'b01111; w[83][191] = 5'b01111; w[83][192] = 5'b01111; w[83][193] = 5'b01111; w[83][194] = 5'b01111; w[83][195] = 5'b01111; w[83][196] = 5'b01111; w[83][197] = 5'b01111; w[83][198] = 5'b01111; w[83][199] = 5'b01111; w[83][200] = 5'b01111; w[83][201] = 5'b01111; w[83][202] = 5'b01111; w[83][203] = 5'b01111; w[83][204] = 5'b01111; w[83][205] = 5'b01111; w[83][206] = 5'b01111; w[83][207] = 5'b01111; w[83][208] = 5'b01111; w[83][209] = 5'b01111; 
w[84][0] = 5'b01111; w[84][1] = 5'b01111; w[84][2] = 5'b01111; w[84][3] = 5'b01111; w[84][4] = 5'b01111; w[84][5] = 5'b01111; w[84][6] = 5'b01111; w[84][7] = 5'b01111; w[84][8] = 5'b01111; w[84][9] = 5'b01111; w[84][10] = 5'b01111; w[84][11] = 5'b01111; w[84][12] = 5'b01111; w[84][13] = 5'b01111; w[84][14] = 5'b01111; w[84][15] = 5'b01111; w[84][16] = 5'b01111; w[84][17] = 5'b01111; w[84][18] = 5'b01111; w[84][19] = 5'b01111; w[84][20] = 5'b01111; w[84][21] = 5'b01111; w[84][22] = 5'b01111; w[84][23] = 5'b01111; w[84][24] = 5'b01111; w[84][25] = 5'b01111; w[84][26] = 5'b01111; w[84][27] = 5'b01111; w[84][28] = 5'b01111; w[84][29] = 5'b01111; w[84][30] = 5'b01111; w[84][31] = 5'b00000; w[84][32] = 5'b10000; w[84][33] = 5'b10000; w[84][34] = 5'b10000; w[84][35] = 5'b10000; w[84][36] = 5'b10000; w[84][37] = 5'b10000; w[84][38] = 5'b00000; w[84][39] = 5'b01111; w[84][40] = 5'b01111; w[84][41] = 5'b01111; w[84][42] = 5'b01111; w[84][43] = 5'b01111; w[84][44] = 5'b01111; w[84][45] = 5'b10000; w[84][46] = 5'b10000; w[84][47] = 5'b10000; w[84][48] = 5'b10000; w[84][49] = 5'b10000; w[84][50] = 5'b10000; w[84][51] = 5'b10000; w[84][52] = 5'b10000; w[84][53] = 5'b01111; w[84][54] = 5'b01111; w[84][55] = 5'b01111; w[84][56] = 5'b01111; w[84][57] = 5'b01111; w[84][58] = 5'b01111; w[84][59] = 5'b00000; w[84][60] = 5'b00000; w[84][61] = 5'b01111; w[84][62] = 5'b10000; w[84][63] = 5'b00000; w[84][64] = 5'b01111; w[84][65] = 5'b00000; w[84][66] = 5'b00000; w[84][67] = 5'b01111; w[84][68] = 5'b01111; w[84][69] = 5'b01111; w[84][70] = 5'b01111; w[84][71] = 5'b01111; w[84][72] = 5'b01111; w[84][73] = 5'b00000; w[84][74] = 5'b01111; w[84][75] = 5'b01111; w[84][76] = 5'b10000; w[84][77] = 5'b00000; w[84][78] = 5'b01111; w[84][79] = 5'b01111; w[84][80] = 5'b00000; w[84][81] = 5'b01111; w[84][82] = 5'b01111; w[84][83] = 5'b01111; w[84][84] = 5'b00000; w[84][85] = 5'b01111; w[84][86] = 5'b01111; w[84][87] = 5'b00000; w[84][88] = 5'b01111; w[84][89] = 5'b01111; w[84][90] = 5'b10000; w[84][91] = 5'b10000; w[84][92] = 5'b01111; w[84][93] = 5'b01111; w[84][94] = 5'b01111; w[84][95] = 5'b01111; w[84][96] = 5'b01111; w[84][97] = 5'b01111; w[84][98] = 5'b01111; w[84][99] = 5'b01111; w[84][100] = 5'b01111; w[84][101] = 5'b00000; w[84][102] = 5'b01111; w[84][103] = 5'b01111; w[84][104] = 5'b10000; w[84][105] = 5'b10000; w[84][106] = 5'b01111; w[84][107] = 5'b00000; w[84][108] = 5'b00000; w[84][109] = 5'b01111; w[84][110] = 5'b01111; w[84][111] = 5'b01111; w[84][112] = 5'b01111; w[84][113] = 5'b01111; w[84][114] = 5'b01111; w[84][115] = 5'b00000; w[84][116] = 5'b01111; w[84][117] = 5'b01111; w[84][118] = 5'b10000; w[84][119] = 5'b10000; w[84][120] = 5'b00000; w[84][121] = 5'b00000; w[84][122] = 5'b00000; w[84][123] = 5'b01111; w[84][124] = 5'b01111; w[84][125] = 5'b01111; w[84][126] = 5'b01111; w[84][127] = 5'b01111; w[84][128] = 5'b01111; w[84][129] = 5'b00000; w[84][130] = 5'b01111; w[84][131] = 5'b01111; w[84][132] = 5'b00000; w[84][133] = 5'b10000; w[84][134] = 5'b01111; w[84][135] = 5'b01111; w[84][136] = 5'b00000; w[84][137] = 5'b01111; w[84][138] = 5'b01111; w[84][139] = 5'b01111; w[84][140] = 5'b01111; w[84][141] = 5'b01111; w[84][142] = 5'b01111; w[84][143] = 5'b00000; w[84][144] = 5'b00000; w[84][145] = 5'b01111; w[84][146] = 5'b00000; w[84][147] = 5'b10000; w[84][148] = 5'b01111; w[84][149] = 5'b00000; w[84][150] = 5'b00000; w[84][151] = 5'b01111; w[84][152] = 5'b01111; w[84][153] = 5'b01111; w[84][154] = 5'b01111; w[84][155] = 5'b01111; w[84][156] = 5'b01111; w[84][157] = 5'b00000; w[84][158] = 5'b00000; w[84][159] = 5'b00000; w[84][160] = 5'b10000; w[84][161] = 5'b10000; w[84][162] = 5'b10000; w[84][163] = 5'b00000; w[84][164] = 5'b00000; w[84][165] = 5'b01111; w[84][166] = 5'b01111; w[84][167] = 5'b01111; w[84][168] = 5'b01111; w[84][169] = 5'b01111; w[84][170] = 5'b01111; w[84][171] = 5'b01111; w[84][172] = 5'b00000; w[84][173] = 5'b00000; w[84][174] = 5'b10000; w[84][175] = 5'b10000; w[84][176] = 5'b10000; w[84][177] = 5'b00000; w[84][178] = 5'b01111; w[84][179] = 5'b01111; w[84][180] = 5'b01111; w[84][181] = 5'b01111; w[84][182] = 5'b01111; w[84][183] = 5'b01111; w[84][184] = 5'b01111; w[84][185] = 5'b01111; w[84][186] = 5'b01111; w[84][187] = 5'b01111; w[84][188] = 5'b01111; w[84][189] = 5'b01111; w[84][190] = 5'b01111; w[84][191] = 5'b01111; w[84][192] = 5'b01111; w[84][193] = 5'b01111; w[84][194] = 5'b01111; w[84][195] = 5'b01111; w[84][196] = 5'b01111; w[84][197] = 5'b01111; w[84][198] = 5'b01111; w[84][199] = 5'b01111; w[84][200] = 5'b01111; w[84][201] = 5'b01111; w[84][202] = 5'b01111; w[84][203] = 5'b01111; w[84][204] = 5'b01111; w[84][205] = 5'b01111; w[84][206] = 5'b01111; w[84][207] = 5'b01111; w[84][208] = 5'b01111; w[84][209] = 5'b01111; 
w[85][0] = 5'b01111; w[85][1] = 5'b01111; w[85][2] = 5'b01111; w[85][3] = 5'b01111; w[85][4] = 5'b01111; w[85][5] = 5'b01111; w[85][6] = 5'b01111; w[85][7] = 5'b01111; w[85][8] = 5'b01111; w[85][9] = 5'b01111; w[85][10] = 5'b01111; w[85][11] = 5'b01111; w[85][12] = 5'b01111; w[85][13] = 5'b01111; w[85][14] = 5'b01111; w[85][15] = 5'b01111; w[85][16] = 5'b01111; w[85][17] = 5'b01111; w[85][18] = 5'b01111; w[85][19] = 5'b01111; w[85][20] = 5'b01111; w[85][21] = 5'b01111; w[85][22] = 5'b01111; w[85][23] = 5'b01111; w[85][24] = 5'b01111; w[85][25] = 5'b01111; w[85][26] = 5'b01111; w[85][27] = 5'b01111; w[85][28] = 5'b01111; w[85][29] = 5'b01111; w[85][30] = 5'b01111; w[85][31] = 5'b00000; w[85][32] = 5'b10000; w[85][33] = 5'b10000; w[85][34] = 5'b10000; w[85][35] = 5'b10000; w[85][36] = 5'b10000; w[85][37] = 5'b10000; w[85][38] = 5'b00000; w[85][39] = 5'b01111; w[85][40] = 5'b01111; w[85][41] = 5'b01111; w[85][42] = 5'b01111; w[85][43] = 5'b01111; w[85][44] = 5'b01111; w[85][45] = 5'b10000; w[85][46] = 5'b10000; w[85][47] = 5'b10000; w[85][48] = 5'b10000; w[85][49] = 5'b10000; w[85][50] = 5'b10000; w[85][51] = 5'b10000; w[85][52] = 5'b10000; w[85][53] = 5'b01111; w[85][54] = 5'b01111; w[85][55] = 5'b01111; w[85][56] = 5'b01111; w[85][57] = 5'b01111; w[85][58] = 5'b01111; w[85][59] = 5'b00000; w[85][60] = 5'b00000; w[85][61] = 5'b01111; w[85][62] = 5'b10000; w[85][63] = 5'b00000; w[85][64] = 5'b01111; w[85][65] = 5'b00000; w[85][66] = 5'b00000; w[85][67] = 5'b01111; w[85][68] = 5'b01111; w[85][69] = 5'b01111; w[85][70] = 5'b01111; w[85][71] = 5'b01111; w[85][72] = 5'b01111; w[85][73] = 5'b00000; w[85][74] = 5'b01111; w[85][75] = 5'b01111; w[85][76] = 5'b10000; w[85][77] = 5'b00000; w[85][78] = 5'b01111; w[85][79] = 5'b01111; w[85][80] = 5'b00000; w[85][81] = 5'b01111; w[85][82] = 5'b01111; w[85][83] = 5'b01111; w[85][84] = 5'b01111; w[85][85] = 5'b00000; w[85][86] = 5'b01111; w[85][87] = 5'b00000; w[85][88] = 5'b01111; w[85][89] = 5'b01111; w[85][90] = 5'b10000; w[85][91] = 5'b10000; w[85][92] = 5'b01111; w[85][93] = 5'b01111; w[85][94] = 5'b01111; w[85][95] = 5'b01111; w[85][96] = 5'b01111; w[85][97] = 5'b01111; w[85][98] = 5'b01111; w[85][99] = 5'b01111; w[85][100] = 5'b01111; w[85][101] = 5'b00000; w[85][102] = 5'b01111; w[85][103] = 5'b01111; w[85][104] = 5'b10000; w[85][105] = 5'b10000; w[85][106] = 5'b01111; w[85][107] = 5'b00000; w[85][108] = 5'b00000; w[85][109] = 5'b01111; w[85][110] = 5'b01111; w[85][111] = 5'b01111; w[85][112] = 5'b01111; w[85][113] = 5'b01111; w[85][114] = 5'b01111; w[85][115] = 5'b00000; w[85][116] = 5'b01111; w[85][117] = 5'b01111; w[85][118] = 5'b10000; w[85][119] = 5'b10000; w[85][120] = 5'b00000; w[85][121] = 5'b00000; w[85][122] = 5'b00000; w[85][123] = 5'b01111; w[85][124] = 5'b01111; w[85][125] = 5'b01111; w[85][126] = 5'b01111; w[85][127] = 5'b01111; w[85][128] = 5'b01111; w[85][129] = 5'b00000; w[85][130] = 5'b01111; w[85][131] = 5'b01111; w[85][132] = 5'b00000; w[85][133] = 5'b10000; w[85][134] = 5'b01111; w[85][135] = 5'b01111; w[85][136] = 5'b00000; w[85][137] = 5'b01111; w[85][138] = 5'b01111; w[85][139] = 5'b01111; w[85][140] = 5'b01111; w[85][141] = 5'b01111; w[85][142] = 5'b01111; w[85][143] = 5'b00000; w[85][144] = 5'b00000; w[85][145] = 5'b01111; w[85][146] = 5'b00000; w[85][147] = 5'b10000; w[85][148] = 5'b01111; w[85][149] = 5'b00000; w[85][150] = 5'b00000; w[85][151] = 5'b01111; w[85][152] = 5'b01111; w[85][153] = 5'b01111; w[85][154] = 5'b01111; w[85][155] = 5'b01111; w[85][156] = 5'b01111; w[85][157] = 5'b00000; w[85][158] = 5'b00000; w[85][159] = 5'b00000; w[85][160] = 5'b10000; w[85][161] = 5'b10000; w[85][162] = 5'b10000; w[85][163] = 5'b00000; w[85][164] = 5'b00000; w[85][165] = 5'b01111; w[85][166] = 5'b01111; w[85][167] = 5'b01111; w[85][168] = 5'b01111; w[85][169] = 5'b01111; w[85][170] = 5'b01111; w[85][171] = 5'b01111; w[85][172] = 5'b00000; w[85][173] = 5'b00000; w[85][174] = 5'b10000; w[85][175] = 5'b10000; w[85][176] = 5'b10000; w[85][177] = 5'b00000; w[85][178] = 5'b01111; w[85][179] = 5'b01111; w[85][180] = 5'b01111; w[85][181] = 5'b01111; w[85][182] = 5'b01111; w[85][183] = 5'b01111; w[85][184] = 5'b01111; w[85][185] = 5'b01111; w[85][186] = 5'b01111; w[85][187] = 5'b01111; w[85][188] = 5'b01111; w[85][189] = 5'b01111; w[85][190] = 5'b01111; w[85][191] = 5'b01111; w[85][192] = 5'b01111; w[85][193] = 5'b01111; w[85][194] = 5'b01111; w[85][195] = 5'b01111; w[85][196] = 5'b01111; w[85][197] = 5'b01111; w[85][198] = 5'b01111; w[85][199] = 5'b01111; w[85][200] = 5'b01111; w[85][201] = 5'b01111; w[85][202] = 5'b01111; w[85][203] = 5'b01111; w[85][204] = 5'b01111; w[85][205] = 5'b01111; w[85][206] = 5'b01111; w[85][207] = 5'b01111; w[85][208] = 5'b01111; w[85][209] = 5'b01111; 
w[86][0] = 5'b01111; w[86][1] = 5'b01111; w[86][2] = 5'b01111; w[86][3] = 5'b01111; w[86][4] = 5'b01111; w[86][5] = 5'b01111; w[86][6] = 5'b01111; w[86][7] = 5'b01111; w[86][8] = 5'b01111; w[86][9] = 5'b01111; w[86][10] = 5'b01111; w[86][11] = 5'b01111; w[86][12] = 5'b01111; w[86][13] = 5'b01111; w[86][14] = 5'b01111; w[86][15] = 5'b01111; w[86][16] = 5'b01111; w[86][17] = 5'b01111; w[86][18] = 5'b01111; w[86][19] = 5'b01111; w[86][20] = 5'b01111; w[86][21] = 5'b01111; w[86][22] = 5'b01111; w[86][23] = 5'b01111; w[86][24] = 5'b01111; w[86][25] = 5'b01111; w[86][26] = 5'b01111; w[86][27] = 5'b01111; w[86][28] = 5'b01111; w[86][29] = 5'b01111; w[86][30] = 5'b00000; w[86][31] = 5'b10000; w[86][32] = 5'b00000; w[86][33] = 5'b10000; w[86][34] = 5'b00000; w[86][35] = 5'b00000; w[86][36] = 5'b00000; w[86][37] = 5'b00000; w[86][38] = 5'b10000; w[86][39] = 5'b00000; w[86][40] = 5'b01111; w[86][41] = 5'b01111; w[86][42] = 5'b01111; w[86][43] = 5'b01111; w[86][44] = 5'b00000; w[86][45] = 5'b00000; w[86][46] = 5'b00000; w[86][47] = 5'b10000; w[86][48] = 5'b00000; w[86][49] = 5'b00000; w[86][50] = 5'b00000; w[86][51] = 5'b00000; w[86][52] = 5'b00000; w[86][53] = 5'b00000; w[86][54] = 5'b01111; w[86][55] = 5'b01111; w[86][56] = 5'b01111; w[86][57] = 5'b01111; w[86][58] = 5'b01111; w[86][59] = 5'b01111; w[86][60] = 5'b01111; w[86][61] = 5'b00000; w[86][62] = 5'b10000; w[86][63] = 5'b10000; w[86][64] = 5'b01111; w[86][65] = 5'b01111; w[86][66] = 5'b01111; w[86][67] = 5'b01111; w[86][68] = 5'b01111; w[86][69] = 5'b01111; w[86][70] = 5'b01111; w[86][71] = 5'b01111; w[86][72] = 5'b01111; w[86][73] = 5'b01111; w[86][74] = 5'b00000; w[86][75] = 5'b00000; w[86][76] = 5'b10000; w[86][77] = 5'b10000; w[86][78] = 5'b01111; w[86][79] = 5'b00000; w[86][80] = 5'b01111; w[86][81] = 5'b01111; w[86][82] = 5'b01111; w[86][83] = 5'b01111; w[86][84] = 5'b01111; w[86][85] = 5'b01111; w[86][86] = 5'b00000; w[86][87] = 5'b01111; w[86][88] = 5'b00000; w[86][89] = 5'b00000; w[86][90] = 5'b10000; w[86][91] = 5'b10000; w[86][92] = 5'b01111; w[86][93] = 5'b00000; w[86][94] = 5'b00000; w[86][95] = 5'b01111; w[86][96] = 5'b01111; w[86][97] = 5'b01111; w[86][98] = 5'b01111; w[86][99] = 5'b01111; w[86][100] = 5'b01111; w[86][101] = 5'b01111; w[86][102] = 5'b00000; w[86][103] = 5'b01111; w[86][104] = 5'b10000; w[86][105] = 5'b10000; w[86][106] = 5'b01111; w[86][107] = 5'b01111; w[86][108] = 5'b01111; w[86][109] = 5'b01111; w[86][110] = 5'b01111; w[86][111] = 5'b01111; w[86][112] = 5'b01111; w[86][113] = 5'b01111; w[86][114] = 5'b01111; w[86][115] = 5'b01111; w[86][116] = 5'b00000; w[86][117] = 5'b01111; w[86][118] = 5'b10000; w[86][119] = 5'b10000; w[86][120] = 5'b01111; w[86][121] = 5'b01111; w[86][122] = 5'b01111; w[86][123] = 5'b01111; w[86][124] = 5'b01111; w[86][125] = 5'b01111; w[86][126] = 5'b01111; w[86][127] = 5'b01111; w[86][128] = 5'b01111; w[86][129] = 5'b01111; w[86][130] = 5'b00000; w[86][131] = 5'b01111; w[86][132] = 5'b10000; w[86][133] = 5'b10000; w[86][134] = 5'b00000; w[86][135] = 5'b00000; w[86][136] = 5'b01111; w[86][137] = 5'b01111; w[86][138] = 5'b01111; w[86][139] = 5'b01111; w[86][140] = 5'b01111; w[86][141] = 5'b01111; w[86][142] = 5'b01111; w[86][143] = 5'b01111; w[86][144] = 5'b01111; w[86][145] = 5'b01111; w[86][146] = 5'b10000; w[86][147] = 5'b10000; w[86][148] = 5'b00000; w[86][149] = 5'b01111; w[86][150] = 5'b01111; w[86][151] = 5'b01111; w[86][152] = 5'b01111; w[86][153] = 5'b01111; w[86][154] = 5'b01111; w[86][155] = 5'b01111; w[86][156] = 5'b01111; w[86][157] = 5'b01111; w[86][158] = 5'b01111; w[86][159] = 5'b01111; w[86][160] = 5'b00000; w[86][161] = 5'b00000; w[86][162] = 5'b00000; w[86][163] = 5'b01111; w[86][164] = 5'b01111; w[86][165] = 5'b01111; w[86][166] = 5'b01111; w[86][167] = 5'b01111; w[86][168] = 5'b01111; w[86][169] = 5'b01111; w[86][170] = 5'b01111; w[86][171] = 5'b00000; w[86][172] = 5'b01111; w[86][173] = 5'b01111; w[86][174] = 5'b00000; w[86][175] = 5'b00000; w[86][176] = 5'b00000; w[86][177] = 5'b01111; w[86][178] = 5'b00000; w[86][179] = 5'b01111; w[86][180] = 5'b01111; w[86][181] = 5'b01111; w[86][182] = 5'b01111; w[86][183] = 5'b01111; w[86][184] = 5'b01111; w[86][185] = 5'b01111; w[86][186] = 5'b01111; w[86][187] = 5'b01111; w[86][188] = 5'b01111; w[86][189] = 5'b01111; w[86][190] = 5'b01111; w[86][191] = 5'b01111; w[86][192] = 5'b01111; w[86][193] = 5'b01111; w[86][194] = 5'b01111; w[86][195] = 5'b01111; w[86][196] = 5'b01111; w[86][197] = 5'b01111; w[86][198] = 5'b01111; w[86][199] = 5'b01111; w[86][200] = 5'b01111; w[86][201] = 5'b01111; w[86][202] = 5'b01111; w[86][203] = 5'b01111; w[86][204] = 5'b01111; w[86][205] = 5'b01111; w[86][206] = 5'b01111; w[86][207] = 5'b01111; w[86][208] = 5'b01111; w[86][209] = 5'b01111; 
w[87][0] = 5'b00000; w[87][1] = 5'b00000; w[87][2] = 5'b00000; w[87][3] = 5'b00000; w[87][4] = 5'b00000; w[87][5] = 5'b00000; w[87][6] = 5'b00000; w[87][7] = 5'b00000; w[87][8] = 5'b00000; w[87][9] = 5'b00000; w[87][10] = 5'b00000; w[87][11] = 5'b00000; w[87][12] = 5'b00000; w[87][13] = 5'b00000; w[87][14] = 5'b00000; w[87][15] = 5'b00000; w[87][16] = 5'b00000; w[87][17] = 5'b00000; w[87][18] = 5'b00000; w[87][19] = 5'b00000; w[87][20] = 5'b00000; w[87][21] = 5'b00000; w[87][22] = 5'b00000; w[87][23] = 5'b00000; w[87][24] = 5'b00000; w[87][25] = 5'b00000; w[87][26] = 5'b00000; w[87][27] = 5'b00000; w[87][28] = 5'b00000; w[87][29] = 5'b00000; w[87][30] = 5'b10000; w[87][31] = 5'b00000; w[87][32] = 5'b01111; w[87][33] = 5'b00000; w[87][34] = 5'b10000; w[87][35] = 5'b10000; w[87][36] = 5'b10000; w[87][37] = 5'b01111; w[87][38] = 5'b00000; w[87][39] = 5'b10000; w[87][40] = 5'b00000; w[87][41] = 5'b00000; w[87][42] = 5'b00000; w[87][43] = 5'b00000; w[87][44] = 5'b10000; w[87][45] = 5'b01111; w[87][46] = 5'b01111; w[87][47] = 5'b00000; w[87][48] = 5'b10000; w[87][49] = 5'b10000; w[87][50] = 5'b10000; w[87][51] = 5'b01111; w[87][52] = 5'b01111; w[87][53] = 5'b10000; w[87][54] = 5'b00000; w[87][55] = 5'b00000; w[87][56] = 5'b00000; w[87][57] = 5'b00000; w[87][58] = 5'b01111; w[87][59] = 5'b01111; w[87][60] = 5'b01111; w[87][61] = 5'b01111; w[87][62] = 5'b10000; w[87][63] = 5'b10000; w[87][64] = 5'b00000; w[87][65] = 5'b01111; w[87][66] = 5'b01111; w[87][67] = 5'b01111; w[87][68] = 5'b00000; w[87][69] = 5'b00000; w[87][70] = 5'b00000; w[87][71] = 5'b00000; w[87][72] = 5'b01111; w[87][73] = 5'b01111; w[87][74] = 5'b01111; w[87][75] = 5'b01111; w[87][76] = 5'b10000; w[87][77] = 5'b10000; w[87][78] = 5'b00000; w[87][79] = 5'b01111; w[87][80] = 5'b01111; w[87][81] = 5'b01111; w[87][82] = 5'b00000; w[87][83] = 5'b00000; w[87][84] = 5'b00000; w[87][85] = 5'b00000; w[87][86] = 5'b01111; w[87][87] = 5'b00000; w[87][88] = 5'b01111; w[87][89] = 5'b01111; w[87][90] = 5'b10000; w[87][91] = 5'b10000; w[87][92] = 5'b00000; w[87][93] = 5'b01111; w[87][94] = 5'b01111; w[87][95] = 5'b00000; w[87][96] = 5'b00000; w[87][97] = 5'b00000; w[87][98] = 5'b00000; w[87][99] = 5'b00000; w[87][100] = 5'b01111; w[87][101] = 5'b01111; w[87][102] = 5'b01111; w[87][103] = 5'b00000; w[87][104] = 5'b10000; w[87][105] = 5'b10000; w[87][106] = 5'b01111; w[87][107] = 5'b01111; w[87][108] = 5'b01111; w[87][109] = 5'b01111; w[87][110] = 5'b00000; w[87][111] = 5'b00000; w[87][112] = 5'b00000; w[87][113] = 5'b00000; w[87][114] = 5'b01111; w[87][115] = 5'b01111; w[87][116] = 5'b01111; w[87][117] = 5'b00000; w[87][118] = 5'b10000; w[87][119] = 5'b10000; w[87][120] = 5'b01111; w[87][121] = 5'b01111; w[87][122] = 5'b01111; w[87][123] = 5'b01111; w[87][124] = 5'b00000; w[87][125] = 5'b00000; w[87][126] = 5'b00000; w[87][127] = 5'b00000; w[87][128] = 5'b01111; w[87][129] = 5'b01111; w[87][130] = 5'b01111; w[87][131] = 5'b00000; w[87][132] = 5'b10000; w[87][133] = 5'b10000; w[87][134] = 5'b01111; w[87][135] = 5'b01111; w[87][136] = 5'b01111; w[87][137] = 5'b01111; w[87][138] = 5'b00000; w[87][139] = 5'b00000; w[87][140] = 5'b00000; w[87][141] = 5'b00000; w[87][142] = 5'b01111; w[87][143] = 5'b01111; w[87][144] = 5'b01111; w[87][145] = 5'b00000; w[87][146] = 5'b10000; w[87][147] = 5'b10000; w[87][148] = 5'b01111; w[87][149] = 5'b01111; w[87][150] = 5'b01111; w[87][151] = 5'b01111; w[87][152] = 5'b00000; w[87][153] = 5'b00000; w[87][154] = 5'b00000; w[87][155] = 5'b00000; w[87][156] = 5'b00000; w[87][157] = 5'b01111; w[87][158] = 5'b01111; w[87][159] = 5'b00000; w[87][160] = 5'b10000; w[87][161] = 5'b10000; w[87][162] = 5'b01111; w[87][163] = 5'b01111; w[87][164] = 5'b01111; w[87][165] = 5'b00000; w[87][166] = 5'b00000; w[87][167] = 5'b00000; w[87][168] = 5'b00000; w[87][169] = 5'b00000; w[87][170] = 5'b00000; w[87][171] = 5'b01111; w[87][172] = 5'b01111; w[87][173] = 5'b00000; w[87][174] = 5'b10000; w[87][175] = 5'b10000; w[87][176] = 5'b01111; w[87][177] = 5'b01111; w[87][178] = 5'b01111; w[87][179] = 5'b00000; w[87][180] = 5'b00000; w[87][181] = 5'b00000; w[87][182] = 5'b00000; w[87][183] = 5'b00000; w[87][184] = 5'b00000; w[87][185] = 5'b00000; w[87][186] = 5'b00000; w[87][187] = 5'b00000; w[87][188] = 5'b00000; w[87][189] = 5'b00000; w[87][190] = 5'b00000; w[87][191] = 5'b00000; w[87][192] = 5'b00000; w[87][193] = 5'b00000; w[87][194] = 5'b00000; w[87][195] = 5'b00000; w[87][196] = 5'b00000; w[87][197] = 5'b00000; w[87][198] = 5'b00000; w[87][199] = 5'b00000; w[87][200] = 5'b00000; w[87][201] = 5'b00000; w[87][202] = 5'b00000; w[87][203] = 5'b00000; w[87][204] = 5'b00000; w[87][205] = 5'b00000; w[87][206] = 5'b00000; w[87][207] = 5'b00000; w[87][208] = 5'b00000; w[87][209] = 5'b00000; 
w[88][0] = 5'b01111; w[88][1] = 5'b01111; w[88][2] = 5'b01111; w[88][3] = 5'b01111; w[88][4] = 5'b01111; w[88][5] = 5'b01111; w[88][6] = 5'b01111; w[88][7] = 5'b01111; w[88][8] = 5'b01111; w[88][9] = 5'b01111; w[88][10] = 5'b01111; w[88][11] = 5'b01111; w[88][12] = 5'b01111; w[88][13] = 5'b01111; w[88][14] = 5'b01111; w[88][15] = 5'b01111; w[88][16] = 5'b01111; w[88][17] = 5'b01111; w[88][18] = 5'b01111; w[88][19] = 5'b01111; w[88][20] = 5'b01111; w[88][21] = 5'b01111; w[88][22] = 5'b01111; w[88][23] = 5'b01111; w[88][24] = 5'b01111; w[88][25] = 5'b01111; w[88][26] = 5'b01111; w[88][27] = 5'b01111; w[88][28] = 5'b01111; w[88][29] = 5'b01111; w[88][30] = 5'b00000; w[88][31] = 5'b01111; w[88][32] = 5'b00000; w[88][33] = 5'b10000; w[88][34] = 5'b10000; w[88][35] = 5'b10000; w[88][36] = 5'b10000; w[88][37] = 5'b00000; w[88][38] = 5'b01111; w[88][39] = 5'b00000; w[88][40] = 5'b01111; w[88][41] = 5'b01111; w[88][42] = 5'b01111; w[88][43] = 5'b01111; w[88][44] = 5'b00000; w[88][45] = 5'b00000; w[88][46] = 5'b00000; w[88][47] = 5'b10000; w[88][48] = 5'b10000; w[88][49] = 5'b10000; w[88][50] = 5'b10000; w[88][51] = 5'b00000; w[88][52] = 5'b00000; w[88][53] = 5'b00000; w[88][54] = 5'b01111; w[88][55] = 5'b01111; w[88][56] = 5'b01111; w[88][57] = 5'b01111; w[88][58] = 5'b00000; w[88][59] = 5'b01111; w[88][60] = 5'b01111; w[88][61] = 5'b01111; w[88][62] = 5'b00000; w[88][63] = 5'b10000; w[88][64] = 5'b01111; w[88][65] = 5'b01111; w[88][66] = 5'b01111; w[88][67] = 5'b00000; w[88][68] = 5'b01111; w[88][69] = 5'b01111; w[88][70] = 5'b01111; w[88][71] = 5'b01111; w[88][72] = 5'b00000; w[88][73] = 5'b01111; w[88][74] = 5'b01111; w[88][75] = 5'b01111; w[88][76] = 5'b00000; w[88][77] = 5'b10000; w[88][78] = 5'b01111; w[88][79] = 5'b01111; w[88][80] = 5'b01111; w[88][81] = 5'b00000; w[88][82] = 5'b01111; w[88][83] = 5'b01111; w[88][84] = 5'b01111; w[88][85] = 5'b01111; w[88][86] = 5'b00000; w[88][87] = 5'b01111; w[88][88] = 5'b00000; w[88][89] = 5'b01111; w[88][90] = 5'b00000; w[88][91] = 5'b00000; w[88][92] = 5'b01111; w[88][93] = 5'b01111; w[88][94] = 5'b01111; w[88][95] = 5'b01111; w[88][96] = 5'b01111; w[88][97] = 5'b01111; w[88][98] = 5'b01111; w[88][99] = 5'b01111; w[88][100] = 5'b00000; w[88][101] = 5'b01111; w[88][102] = 5'b01111; w[88][103] = 5'b01111; w[88][104] = 5'b00000; w[88][105] = 5'b00000; w[88][106] = 5'b00000; w[88][107] = 5'b01111; w[88][108] = 5'b01111; w[88][109] = 5'b00000; w[88][110] = 5'b01111; w[88][111] = 5'b01111; w[88][112] = 5'b01111; w[88][113] = 5'b01111; w[88][114] = 5'b00000; w[88][115] = 5'b01111; w[88][116] = 5'b01111; w[88][117] = 5'b01111; w[88][118] = 5'b00000; w[88][119] = 5'b00000; w[88][120] = 5'b01111; w[88][121] = 5'b01111; w[88][122] = 5'b01111; w[88][123] = 5'b00000; w[88][124] = 5'b01111; w[88][125] = 5'b01111; w[88][126] = 5'b01111; w[88][127] = 5'b01111; w[88][128] = 5'b00000; w[88][129] = 5'b01111; w[88][130] = 5'b01111; w[88][131] = 5'b01111; w[88][132] = 5'b10000; w[88][133] = 5'b00000; w[88][134] = 5'b01111; w[88][135] = 5'b01111; w[88][136] = 5'b01111; w[88][137] = 5'b00000; w[88][138] = 5'b01111; w[88][139] = 5'b01111; w[88][140] = 5'b01111; w[88][141] = 5'b01111; w[88][142] = 5'b00000; w[88][143] = 5'b01111; w[88][144] = 5'b01111; w[88][145] = 5'b01111; w[88][146] = 5'b10000; w[88][147] = 5'b00000; w[88][148] = 5'b01111; w[88][149] = 5'b01111; w[88][150] = 5'b01111; w[88][151] = 5'b00000; w[88][152] = 5'b01111; w[88][153] = 5'b01111; w[88][154] = 5'b01111; w[88][155] = 5'b01111; w[88][156] = 5'b01111; w[88][157] = 5'b01111; w[88][158] = 5'b01111; w[88][159] = 5'b10000; w[88][160] = 5'b10000; w[88][161] = 5'b10000; w[88][162] = 5'b00000; w[88][163] = 5'b01111; w[88][164] = 5'b01111; w[88][165] = 5'b01111; w[88][166] = 5'b01111; w[88][167] = 5'b01111; w[88][168] = 5'b01111; w[88][169] = 5'b01111; w[88][170] = 5'b01111; w[88][171] = 5'b01111; w[88][172] = 5'b01111; w[88][173] = 5'b10000; w[88][174] = 5'b10000; w[88][175] = 5'b10000; w[88][176] = 5'b00000; w[88][177] = 5'b01111; w[88][178] = 5'b01111; w[88][179] = 5'b01111; w[88][180] = 5'b01111; w[88][181] = 5'b01111; w[88][182] = 5'b01111; w[88][183] = 5'b01111; w[88][184] = 5'b01111; w[88][185] = 5'b01111; w[88][186] = 5'b01111; w[88][187] = 5'b01111; w[88][188] = 5'b01111; w[88][189] = 5'b01111; w[88][190] = 5'b01111; w[88][191] = 5'b01111; w[88][192] = 5'b01111; w[88][193] = 5'b01111; w[88][194] = 5'b01111; w[88][195] = 5'b01111; w[88][196] = 5'b01111; w[88][197] = 5'b01111; w[88][198] = 5'b01111; w[88][199] = 5'b01111; w[88][200] = 5'b01111; w[88][201] = 5'b01111; w[88][202] = 5'b01111; w[88][203] = 5'b01111; w[88][204] = 5'b01111; w[88][205] = 5'b01111; w[88][206] = 5'b01111; w[88][207] = 5'b01111; w[88][208] = 5'b01111; w[88][209] = 5'b01111; 
w[89][0] = 5'b01111; w[89][1] = 5'b01111; w[89][2] = 5'b01111; w[89][3] = 5'b01111; w[89][4] = 5'b01111; w[89][5] = 5'b01111; w[89][6] = 5'b01111; w[89][7] = 5'b01111; w[89][8] = 5'b01111; w[89][9] = 5'b01111; w[89][10] = 5'b01111; w[89][11] = 5'b01111; w[89][12] = 5'b01111; w[89][13] = 5'b01111; w[89][14] = 5'b01111; w[89][15] = 5'b01111; w[89][16] = 5'b01111; w[89][17] = 5'b01111; w[89][18] = 5'b01111; w[89][19] = 5'b01111; w[89][20] = 5'b01111; w[89][21] = 5'b01111; w[89][22] = 5'b01111; w[89][23] = 5'b01111; w[89][24] = 5'b01111; w[89][25] = 5'b01111; w[89][26] = 5'b01111; w[89][27] = 5'b01111; w[89][28] = 5'b01111; w[89][29] = 5'b01111; w[89][30] = 5'b00000; w[89][31] = 5'b01111; w[89][32] = 5'b00000; w[89][33] = 5'b10000; w[89][34] = 5'b10000; w[89][35] = 5'b10000; w[89][36] = 5'b10000; w[89][37] = 5'b00000; w[89][38] = 5'b01111; w[89][39] = 5'b00000; w[89][40] = 5'b01111; w[89][41] = 5'b01111; w[89][42] = 5'b01111; w[89][43] = 5'b01111; w[89][44] = 5'b00000; w[89][45] = 5'b00000; w[89][46] = 5'b00000; w[89][47] = 5'b10000; w[89][48] = 5'b10000; w[89][49] = 5'b10000; w[89][50] = 5'b10000; w[89][51] = 5'b00000; w[89][52] = 5'b00000; w[89][53] = 5'b00000; w[89][54] = 5'b01111; w[89][55] = 5'b01111; w[89][56] = 5'b01111; w[89][57] = 5'b01111; w[89][58] = 5'b00000; w[89][59] = 5'b01111; w[89][60] = 5'b01111; w[89][61] = 5'b01111; w[89][62] = 5'b00000; w[89][63] = 5'b10000; w[89][64] = 5'b01111; w[89][65] = 5'b01111; w[89][66] = 5'b01111; w[89][67] = 5'b00000; w[89][68] = 5'b01111; w[89][69] = 5'b01111; w[89][70] = 5'b01111; w[89][71] = 5'b01111; w[89][72] = 5'b00000; w[89][73] = 5'b01111; w[89][74] = 5'b01111; w[89][75] = 5'b01111; w[89][76] = 5'b00000; w[89][77] = 5'b10000; w[89][78] = 5'b01111; w[89][79] = 5'b01111; w[89][80] = 5'b01111; w[89][81] = 5'b00000; w[89][82] = 5'b01111; w[89][83] = 5'b01111; w[89][84] = 5'b01111; w[89][85] = 5'b01111; w[89][86] = 5'b00000; w[89][87] = 5'b01111; w[89][88] = 5'b01111; w[89][89] = 5'b00000; w[89][90] = 5'b00000; w[89][91] = 5'b00000; w[89][92] = 5'b01111; w[89][93] = 5'b01111; w[89][94] = 5'b01111; w[89][95] = 5'b01111; w[89][96] = 5'b01111; w[89][97] = 5'b01111; w[89][98] = 5'b01111; w[89][99] = 5'b01111; w[89][100] = 5'b00000; w[89][101] = 5'b01111; w[89][102] = 5'b01111; w[89][103] = 5'b01111; w[89][104] = 5'b00000; w[89][105] = 5'b00000; w[89][106] = 5'b00000; w[89][107] = 5'b01111; w[89][108] = 5'b01111; w[89][109] = 5'b00000; w[89][110] = 5'b01111; w[89][111] = 5'b01111; w[89][112] = 5'b01111; w[89][113] = 5'b01111; w[89][114] = 5'b00000; w[89][115] = 5'b01111; w[89][116] = 5'b01111; w[89][117] = 5'b01111; w[89][118] = 5'b00000; w[89][119] = 5'b00000; w[89][120] = 5'b01111; w[89][121] = 5'b01111; w[89][122] = 5'b01111; w[89][123] = 5'b00000; w[89][124] = 5'b01111; w[89][125] = 5'b01111; w[89][126] = 5'b01111; w[89][127] = 5'b01111; w[89][128] = 5'b00000; w[89][129] = 5'b01111; w[89][130] = 5'b01111; w[89][131] = 5'b01111; w[89][132] = 5'b10000; w[89][133] = 5'b00000; w[89][134] = 5'b01111; w[89][135] = 5'b01111; w[89][136] = 5'b01111; w[89][137] = 5'b00000; w[89][138] = 5'b01111; w[89][139] = 5'b01111; w[89][140] = 5'b01111; w[89][141] = 5'b01111; w[89][142] = 5'b00000; w[89][143] = 5'b01111; w[89][144] = 5'b01111; w[89][145] = 5'b01111; w[89][146] = 5'b10000; w[89][147] = 5'b00000; w[89][148] = 5'b01111; w[89][149] = 5'b01111; w[89][150] = 5'b01111; w[89][151] = 5'b00000; w[89][152] = 5'b01111; w[89][153] = 5'b01111; w[89][154] = 5'b01111; w[89][155] = 5'b01111; w[89][156] = 5'b01111; w[89][157] = 5'b01111; w[89][158] = 5'b01111; w[89][159] = 5'b10000; w[89][160] = 5'b10000; w[89][161] = 5'b10000; w[89][162] = 5'b00000; w[89][163] = 5'b01111; w[89][164] = 5'b01111; w[89][165] = 5'b01111; w[89][166] = 5'b01111; w[89][167] = 5'b01111; w[89][168] = 5'b01111; w[89][169] = 5'b01111; w[89][170] = 5'b01111; w[89][171] = 5'b01111; w[89][172] = 5'b01111; w[89][173] = 5'b10000; w[89][174] = 5'b10000; w[89][175] = 5'b10000; w[89][176] = 5'b00000; w[89][177] = 5'b01111; w[89][178] = 5'b01111; w[89][179] = 5'b01111; w[89][180] = 5'b01111; w[89][181] = 5'b01111; w[89][182] = 5'b01111; w[89][183] = 5'b01111; w[89][184] = 5'b01111; w[89][185] = 5'b01111; w[89][186] = 5'b01111; w[89][187] = 5'b01111; w[89][188] = 5'b01111; w[89][189] = 5'b01111; w[89][190] = 5'b01111; w[89][191] = 5'b01111; w[89][192] = 5'b01111; w[89][193] = 5'b01111; w[89][194] = 5'b01111; w[89][195] = 5'b01111; w[89][196] = 5'b01111; w[89][197] = 5'b01111; w[89][198] = 5'b01111; w[89][199] = 5'b01111; w[89][200] = 5'b01111; w[89][201] = 5'b01111; w[89][202] = 5'b01111; w[89][203] = 5'b01111; w[89][204] = 5'b01111; w[89][205] = 5'b01111; w[89][206] = 5'b01111; w[89][207] = 5'b01111; w[89][208] = 5'b01111; w[89][209] = 5'b01111; 
w[90][0] = 5'b10000; w[90][1] = 5'b10000; w[90][2] = 5'b10000; w[90][3] = 5'b10000; w[90][4] = 5'b10000; w[90][5] = 5'b10000; w[90][6] = 5'b10000; w[90][7] = 5'b10000; w[90][8] = 5'b10000; w[90][9] = 5'b10000; w[90][10] = 5'b10000; w[90][11] = 5'b10000; w[90][12] = 5'b10000; w[90][13] = 5'b10000; w[90][14] = 5'b10000; w[90][15] = 5'b10000; w[90][16] = 5'b10000; w[90][17] = 5'b10000; w[90][18] = 5'b10000; w[90][19] = 5'b10000; w[90][20] = 5'b10000; w[90][21] = 5'b10000; w[90][22] = 5'b10000; w[90][23] = 5'b10000; w[90][24] = 5'b10000; w[90][25] = 5'b10000; w[90][26] = 5'b10000; w[90][27] = 5'b10000; w[90][28] = 5'b10000; w[90][29] = 5'b10000; w[90][30] = 5'b00000; w[90][31] = 5'b01111; w[90][32] = 5'b00000; w[90][33] = 5'b01111; w[90][34] = 5'b00000; w[90][35] = 5'b00000; w[90][36] = 5'b00000; w[90][37] = 5'b00000; w[90][38] = 5'b01111; w[90][39] = 5'b00000; w[90][40] = 5'b10000; w[90][41] = 5'b10000; w[90][42] = 5'b10000; w[90][43] = 5'b10000; w[90][44] = 5'b00000; w[90][45] = 5'b00000; w[90][46] = 5'b00000; w[90][47] = 5'b01111; w[90][48] = 5'b00000; w[90][49] = 5'b00000; w[90][50] = 5'b00000; w[90][51] = 5'b00000; w[90][52] = 5'b00000; w[90][53] = 5'b00000; w[90][54] = 5'b10000; w[90][55] = 5'b10000; w[90][56] = 5'b10000; w[90][57] = 5'b10000; w[90][58] = 5'b10000; w[90][59] = 5'b10000; w[90][60] = 5'b10000; w[90][61] = 5'b00000; w[90][62] = 5'b01111; w[90][63] = 5'b01111; w[90][64] = 5'b10000; w[90][65] = 5'b10000; w[90][66] = 5'b10000; w[90][67] = 5'b10000; w[90][68] = 5'b10000; w[90][69] = 5'b10000; w[90][70] = 5'b10000; w[90][71] = 5'b10000; w[90][72] = 5'b10000; w[90][73] = 5'b10000; w[90][74] = 5'b00000; w[90][75] = 5'b00000; w[90][76] = 5'b01111; w[90][77] = 5'b01111; w[90][78] = 5'b10000; w[90][79] = 5'b00000; w[90][80] = 5'b10000; w[90][81] = 5'b10000; w[90][82] = 5'b10000; w[90][83] = 5'b10000; w[90][84] = 5'b10000; w[90][85] = 5'b10000; w[90][86] = 5'b10000; w[90][87] = 5'b10000; w[90][88] = 5'b00000; w[90][89] = 5'b00000; w[90][90] = 5'b00000; w[90][91] = 5'b01111; w[90][92] = 5'b10000; w[90][93] = 5'b00000; w[90][94] = 5'b00000; w[90][95] = 5'b10000; w[90][96] = 5'b10000; w[90][97] = 5'b10000; w[90][98] = 5'b10000; w[90][99] = 5'b10000; w[90][100] = 5'b10000; w[90][101] = 5'b10000; w[90][102] = 5'b00000; w[90][103] = 5'b10000; w[90][104] = 5'b01111; w[90][105] = 5'b01111; w[90][106] = 5'b10000; w[90][107] = 5'b10000; w[90][108] = 5'b10000; w[90][109] = 5'b10000; w[90][110] = 5'b10000; w[90][111] = 5'b10000; w[90][112] = 5'b10000; w[90][113] = 5'b10000; w[90][114] = 5'b10000; w[90][115] = 5'b10000; w[90][116] = 5'b00000; w[90][117] = 5'b10000; w[90][118] = 5'b01111; w[90][119] = 5'b01111; w[90][120] = 5'b10000; w[90][121] = 5'b10000; w[90][122] = 5'b10000; w[90][123] = 5'b10000; w[90][124] = 5'b10000; w[90][125] = 5'b10000; w[90][126] = 5'b10000; w[90][127] = 5'b10000; w[90][128] = 5'b10000; w[90][129] = 5'b10000; w[90][130] = 5'b00000; w[90][131] = 5'b10000; w[90][132] = 5'b01111; w[90][133] = 5'b01111; w[90][134] = 5'b00000; w[90][135] = 5'b00000; w[90][136] = 5'b10000; w[90][137] = 5'b10000; w[90][138] = 5'b10000; w[90][139] = 5'b10000; w[90][140] = 5'b10000; w[90][141] = 5'b10000; w[90][142] = 5'b10000; w[90][143] = 5'b10000; w[90][144] = 5'b10000; w[90][145] = 5'b10000; w[90][146] = 5'b01111; w[90][147] = 5'b01111; w[90][148] = 5'b00000; w[90][149] = 5'b10000; w[90][150] = 5'b10000; w[90][151] = 5'b10000; w[90][152] = 5'b10000; w[90][153] = 5'b10000; w[90][154] = 5'b10000; w[90][155] = 5'b10000; w[90][156] = 5'b10000; w[90][157] = 5'b10000; w[90][158] = 5'b10000; w[90][159] = 5'b10000; w[90][160] = 5'b00000; w[90][161] = 5'b00000; w[90][162] = 5'b00000; w[90][163] = 5'b10000; w[90][164] = 5'b10000; w[90][165] = 5'b10000; w[90][166] = 5'b10000; w[90][167] = 5'b10000; w[90][168] = 5'b10000; w[90][169] = 5'b10000; w[90][170] = 5'b10000; w[90][171] = 5'b00000; w[90][172] = 5'b10000; w[90][173] = 5'b10000; w[90][174] = 5'b00000; w[90][175] = 5'b00000; w[90][176] = 5'b00000; w[90][177] = 5'b10000; w[90][178] = 5'b00000; w[90][179] = 5'b10000; w[90][180] = 5'b10000; w[90][181] = 5'b10000; w[90][182] = 5'b10000; w[90][183] = 5'b10000; w[90][184] = 5'b10000; w[90][185] = 5'b10000; w[90][186] = 5'b10000; w[90][187] = 5'b10000; w[90][188] = 5'b10000; w[90][189] = 5'b10000; w[90][190] = 5'b10000; w[90][191] = 5'b10000; w[90][192] = 5'b10000; w[90][193] = 5'b10000; w[90][194] = 5'b10000; w[90][195] = 5'b10000; w[90][196] = 5'b10000; w[90][197] = 5'b10000; w[90][198] = 5'b10000; w[90][199] = 5'b10000; w[90][200] = 5'b10000; w[90][201] = 5'b10000; w[90][202] = 5'b10000; w[90][203] = 5'b10000; w[90][204] = 5'b10000; w[90][205] = 5'b10000; w[90][206] = 5'b10000; w[90][207] = 5'b10000; w[90][208] = 5'b10000; w[90][209] = 5'b10000; 
w[91][0] = 5'b10000; w[91][1] = 5'b10000; w[91][2] = 5'b10000; w[91][3] = 5'b10000; w[91][4] = 5'b10000; w[91][5] = 5'b10000; w[91][6] = 5'b10000; w[91][7] = 5'b10000; w[91][8] = 5'b10000; w[91][9] = 5'b10000; w[91][10] = 5'b10000; w[91][11] = 5'b10000; w[91][12] = 5'b10000; w[91][13] = 5'b10000; w[91][14] = 5'b10000; w[91][15] = 5'b10000; w[91][16] = 5'b10000; w[91][17] = 5'b10000; w[91][18] = 5'b10000; w[91][19] = 5'b10000; w[91][20] = 5'b10000; w[91][21] = 5'b10000; w[91][22] = 5'b10000; w[91][23] = 5'b10000; w[91][24] = 5'b10000; w[91][25] = 5'b10000; w[91][26] = 5'b10000; w[91][27] = 5'b10000; w[91][28] = 5'b10000; w[91][29] = 5'b10000; w[91][30] = 5'b00000; w[91][31] = 5'b01111; w[91][32] = 5'b00000; w[91][33] = 5'b01111; w[91][34] = 5'b00000; w[91][35] = 5'b00000; w[91][36] = 5'b00000; w[91][37] = 5'b00000; w[91][38] = 5'b01111; w[91][39] = 5'b00000; w[91][40] = 5'b10000; w[91][41] = 5'b10000; w[91][42] = 5'b10000; w[91][43] = 5'b10000; w[91][44] = 5'b00000; w[91][45] = 5'b00000; w[91][46] = 5'b00000; w[91][47] = 5'b01111; w[91][48] = 5'b00000; w[91][49] = 5'b00000; w[91][50] = 5'b00000; w[91][51] = 5'b00000; w[91][52] = 5'b00000; w[91][53] = 5'b00000; w[91][54] = 5'b10000; w[91][55] = 5'b10000; w[91][56] = 5'b10000; w[91][57] = 5'b10000; w[91][58] = 5'b10000; w[91][59] = 5'b10000; w[91][60] = 5'b10000; w[91][61] = 5'b00000; w[91][62] = 5'b01111; w[91][63] = 5'b01111; w[91][64] = 5'b10000; w[91][65] = 5'b10000; w[91][66] = 5'b10000; w[91][67] = 5'b10000; w[91][68] = 5'b10000; w[91][69] = 5'b10000; w[91][70] = 5'b10000; w[91][71] = 5'b10000; w[91][72] = 5'b10000; w[91][73] = 5'b10000; w[91][74] = 5'b00000; w[91][75] = 5'b00000; w[91][76] = 5'b01111; w[91][77] = 5'b01111; w[91][78] = 5'b10000; w[91][79] = 5'b00000; w[91][80] = 5'b10000; w[91][81] = 5'b10000; w[91][82] = 5'b10000; w[91][83] = 5'b10000; w[91][84] = 5'b10000; w[91][85] = 5'b10000; w[91][86] = 5'b10000; w[91][87] = 5'b10000; w[91][88] = 5'b00000; w[91][89] = 5'b00000; w[91][90] = 5'b01111; w[91][91] = 5'b00000; w[91][92] = 5'b10000; w[91][93] = 5'b00000; w[91][94] = 5'b00000; w[91][95] = 5'b10000; w[91][96] = 5'b10000; w[91][97] = 5'b10000; w[91][98] = 5'b10000; w[91][99] = 5'b10000; w[91][100] = 5'b10000; w[91][101] = 5'b10000; w[91][102] = 5'b00000; w[91][103] = 5'b10000; w[91][104] = 5'b01111; w[91][105] = 5'b01111; w[91][106] = 5'b10000; w[91][107] = 5'b10000; w[91][108] = 5'b10000; w[91][109] = 5'b10000; w[91][110] = 5'b10000; w[91][111] = 5'b10000; w[91][112] = 5'b10000; w[91][113] = 5'b10000; w[91][114] = 5'b10000; w[91][115] = 5'b10000; w[91][116] = 5'b00000; w[91][117] = 5'b10000; w[91][118] = 5'b01111; w[91][119] = 5'b01111; w[91][120] = 5'b10000; w[91][121] = 5'b10000; w[91][122] = 5'b10000; w[91][123] = 5'b10000; w[91][124] = 5'b10000; w[91][125] = 5'b10000; w[91][126] = 5'b10000; w[91][127] = 5'b10000; w[91][128] = 5'b10000; w[91][129] = 5'b10000; w[91][130] = 5'b00000; w[91][131] = 5'b10000; w[91][132] = 5'b01111; w[91][133] = 5'b01111; w[91][134] = 5'b00000; w[91][135] = 5'b00000; w[91][136] = 5'b10000; w[91][137] = 5'b10000; w[91][138] = 5'b10000; w[91][139] = 5'b10000; w[91][140] = 5'b10000; w[91][141] = 5'b10000; w[91][142] = 5'b10000; w[91][143] = 5'b10000; w[91][144] = 5'b10000; w[91][145] = 5'b10000; w[91][146] = 5'b01111; w[91][147] = 5'b01111; w[91][148] = 5'b00000; w[91][149] = 5'b10000; w[91][150] = 5'b10000; w[91][151] = 5'b10000; w[91][152] = 5'b10000; w[91][153] = 5'b10000; w[91][154] = 5'b10000; w[91][155] = 5'b10000; w[91][156] = 5'b10000; w[91][157] = 5'b10000; w[91][158] = 5'b10000; w[91][159] = 5'b10000; w[91][160] = 5'b00000; w[91][161] = 5'b00000; w[91][162] = 5'b00000; w[91][163] = 5'b10000; w[91][164] = 5'b10000; w[91][165] = 5'b10000; w[91][166] = 5'b10000; w[91][167] = 5'b10000; w[91][168] = 5'b10000; w[91][169] = 5'b10000; w[91][170] = 5'b10000; w[91][171] = 5'b00000; w[91][172] = 5'b10000; w[91][173] = 5'b10000; w[91][174] = 5'b00000; w[91][175] = 5'b00000; w[91][176] = 5'b00000; w[91][177] = 5'b10000; w[91][178] = 5'b00000; w[91][179] = 5'b10000; w[91][180] = 5'b10000; w[91][181] = 5'b10000; w[91][182] = 5'b10000; w[91][183] = 5'b10000; w[91][184] = 5'b10000; w[91][185] = 5'b10000; w[91][186] = 5'b10000; w[91][187] = 5'b10000; w[91][188] = 5'b10000; w[91][189] = 5'b10000; w[91][190] = 5'b10000; w[91][191] = 5'b10000; w[91][192] = 5'b10000; w[91][193] = 5'b10000; w[91][194] = 5'b10000; w[91][195] = 5'b10000; w[91][196] = 5'b10000; w[91][197] = 5'b10000; w[91][198] = 5'b10000; w[91][199] = 5'b10000; w[91][200] = 5'b10000; w[91][201] = 5'b10000; w[91][202] = 5'b10000; w[91][203] = 5'b10000; w[91][204] = 5'b10000; w[91][205] = 5'b10000; w[91][206] = 5'b10000; w[91][207] = 5'b10000; w[91][208] = 5'b10000; w[91][209] = 5'b10000; 
w[92][0] = 5'b01111; w[92][1] = 5'b01111; w[92][2] = 5'b01111; w[92][3] = 5'b01111; w[92][4] = 5'b01111; w[92][5] = 5'b01111; w[92][6] = 5'b01111; w[92][7] = 5'b01111; w[92][8] = 5'b01111; w[92][9] = 5'b01111; w[92][10] = 5'b01111; w[92][11] = 5'b01111; w[92][12] = 5'b01111; w[92][13] = 5'b01111; w[92][14] = 5'b01111; w[92][15] = 5'b01111; w[92][16] = 5'b01111; w[92][17] = 5'b01111; w[92][18] = 5'b01111; w[92][19] = 5'b01111; w[92][20] = 5'b01111; w[92][21] = 5'b01111; w[92][22] = 5'b01111; w[92][23] = 5'b01111; w[92][24] = 5'b01111; w[92][25] = 5'b01111; w[92][26] = 5'b01111; w[92][27] = 5'b01111; w[92][28] = 5'b01111; w[92][29] = 5'b01111; w[92][30] = 5'b01111; w[92][31] = 5'b00000; w[92][32] = 5'b10000; w[92][33] = 5'b10000; w[92][34] = 5'b10000; w[92][35] = 5'b10000; w[92][36] = 5'b10000; w[92][37] = 5'b10000; w[92][38] = 5'b00000; w[92][39] = 5'b01111; w[92][40] = 5'b01111; w[92][41] = 5'b01111; w[92][42] = 5'b01111; w[92][43] = 5'b01111; w[92][44] = 5'b01111; w[92][45] = 5'b10000; w[92][46] = 5'b10000; w[92][47] = 5'b10000; w[92][48] = 5'b10000; w[92][49] = 5'b10000; w[92][50] = 5'b10000; w[92][51] = 5'b10000; w[92][52] = 5'b10000; w[92][53] = 5'b01111; w[92][54] = 5'b01111; w[92][55] = 5'b01111; w[92][56] = 5'b01111; w[92][57] = 5'b01111; w[92][58] = 5'b01111; w[92][59] = 5'b00000; w[92][60] = 5'b00000; w[92][61] = 5'b01111; w[92][62] = 5'b10000; w[92][63] = 5'b00000; w[92][64] = 5'b01111; w[92][65] = 5'b00000; w[92][66] = 5'b00000; w[92][67] = 5'b01111; w[92][68] = 5'b01111; w[92][69] = 5'b01111; w[92][70] = 5'b01111; w[92][71] = 5'b01111; w[92][72] = 5'b01111; w[92][73] = 5'b00000; w[92][74] = 5'b01111; w[92][75] = 5'b01111; w[92][76] = 5'b10000; w[92][77] = 5'b00000; w[92][78] = 5'b01111; w[92][79] = 5'b01111; w[92][80] = 5'b00000; w[92][81] = 5'b01111; w[92][82] = 5'b01111; w[92][83] = 5'b01111; w[92][84] = 5'b01111; w[92][85] = 5'b01111; w[92][86] = 5'b01111; w[92][87] = 5'b00000; w[92][88] = 5'b01111; w[92][89] = 5'b01111; w[92][90] = 5'b10000; w[92][91] = 5'b10000; w[92][92] = 5'b00000; w[92][93] = 5'b01111; w[92][94] = 5'b01111; w[92][95] = 5'b01111; w[92][96] = 5'b01111; w[92][97] = 5'b01111; w[92][98] = 5'b01111; w[92][99] = 5'b01111; w[92][100] = 5'b01111; w[92][101] = 5'b00000; w[92][102] = 5'b01111; w[92][103] = 5'b01111; w[92][104] = 5'b10000; w[92][105] = 5'b10000; w[92][106] = 5'b01111; w[92][107] = 5'b00000; w[92][108] = 5'b00000; w[92][109] = 5'b01111; w[92][110] = 5'b01111; w[92][111] = 5'b01111; w[92][112] = 5'b01111; w[92][113] = 5'b01111; w[92][114] = 5'b01111; w[92][115] = 5'b00000; w[92][116] = 5'b01111; w[92][117] = 5'b01111; w[92][118] = 5'b10000; w[92][119] = 5'b10000; w[92][120] = 5'b00000; w[92][121] = 5'b00000; w[92][122] = 5'b00000; w[92][123] = 5'b01111; w[92][124] = 5'b01111; w[92][125] = 5'b01111; w[92][126] = 5'b01111; w[92][127] = 5'b01111; w[92][128] = 5'b01111; w[92][129] = 5'b00000; w[92][130] = 5'b01111; w[92][131] = 5'b01111; w[92][132] = 5'b00000; w[92][133] = 5'b10000; w[92][134] = 5'b01111; w[92][135] = 5'b01111; w[92][136] = 5'b00000; w[92][137] = 5'b01111; w[92][138] = 5'b01111; w[92][139] = 5'b01111; w[92][140] = 5'b01111; w[92][141] = 5'b01111; w[92][142] = 5'b01111; w[92][143] = 5'b00000; w[92][144] = 5'b00000; w[92][145] = 5'b01111; w[92][146] = 5'b00000; w[92][147] = 5'b10000; w[92][148] = 5'b01111; w[92][149] = 5'b00000; w[92][150] = 5'b00000; w[92][151] = 5'b01111; w[92][152] = 5'b01111; w[92][153] = 5'b01111; w[92][154] = 5'b01111; w[92][155] = 5'b01111; w[92][156] = 5'b01111; w[92][157] = 5'b00000; w[92][158] = 5'b00000; w[92][159] = 5'b00000; w[92][160] = 5'b10000; w[92][161] = 5'b10000; w[92][162] = 5'b10000; w[92][163] = 5'b00000; w[92][164] = 5'b00000; w[92][165] = 5'b01111; w[92][166] = 5'b01111; w[92][167] = 5'b01111; w[92][168] = 5'b01111; w[92][169] = 5'b01111; w[92][170] = 5'b01111; w[92][171] = 5'b01111; w[92][172] = 5'b00000; w[92][173] = 5'b00000; w[92][174] = 5'b10000; w[92][175] = 5'b10000; w[92][176] = 5'b10000; w[92][177] = 5'b00000; w[92][178] = 5'b01111; w[92][179] = 5'b01111; w[92][180] = 5'b01111; w[92][181] = 5'b01111; w[92][182] = 5'b01111; w[92][183] = 5'b01111; w[92][184] = 5'b01111; w[92][185] = 5'b01111; w[92][186] = 5'b01111; w[92][187] = 5'b01111; w[92][188] = 5'b01111; w[92][189] = 5'b01111; w[92][190] = 5'b01111; w[92][191] = 5'b01111; w[92][192] = 5'b01111; w[92][193] = 5'b01111; w[92][194] = 5'b01111; w[92][195] = 5'b01111; w[92][196] = 5'b01111; w[92][197] = 5'b01111; w[92][198] = 5'b01111; w[92][199] = 5'b01111; w[92][200] = 5'b01111; w[92][201] = 5'b01111; w[92][202] = 5'b01111; w[92][203] = 5'b01111; w[92][204] = 5'b01111; w[92][205] = 5'b01111; w[92][206] = 5'b01111; w[92][207] = 5'b01111; w[92][208] = 5'b01111; w[92][209] = 5'b01111; 
w[93][0] = 5'b01111; w[93][1] = 5'b01111; w[93][2] = 5'b01111; w[93][3] = 5'b01111; w[93][4] = 5'b01111; w[93][5] = 5'b01111; w[93][6] = 5'b01111; w[93][7] = 5'b01111; w[93][8] = 5'b01111; w[93][9] = 5'b01111; w[93][10] = 5'b01111; w[93][11] = 5'b01111; w[93][12] = 5'b01111; w[93][13] = 5'b01111; w[93][14] = 5'b01111; w[93][15] = 5'b01111; w[93][16] = 5'b01111; w[93][17] = 5'b01111; w[93][18] = 5'b01111; w[93][19] = 5'b01111; w[93][20] = 5'b01111; w[93][21] = 5'b01111; w[93][22] = 5'b01111; w[93][23] = 5'b01111; w[93][24] = 5'b01111; w[93][25] = 5'b01111; w[93][26] = 5'b01111; w[93][27] = 5'b01111; w[93][28] = 5'b01111; w[93][29] = 5'b01111; w[93][30] = 5'b00000; w[93][31] = 5'b01111; w[93][32] = 5'b00000; w[93][33] = 5'b10000; w[93][34] = 5'b10000; w[93][35] = 5'b10000; w[93][36] = 5'b10000; w[93][37] = 5'b00000; w[93][38] = 5'b01111; w[93][39] = 5'b00000; w[93][40] = 5'b01111; w[93][41] = 5'b01111; w[93][42] = 5'b01111; w[93][43] = 5'b01111; w[93][44] = 5'b00000; w[93][45] = 5'b00000; w[93][46] = 5'b00000; w[93][47] = 5'b10000; w[93][48] = 5'b10000; w[93][49] = 5'b10000; w[93][50] = 5'b10000; w[93][51] = 5'b00000; w[93][52] = 5'b00000; w[93][53] = 5'b00000; w[93][54] = 5'b01111; w[93][55] = 5'b01111; w[93][56] = 5'b01111; w[93][57] = 5'b01111; w[93][58] = 5'b00000; w[93][59] = 5'b01111; w[93][60] = 5'b01111; w[93][61] = 5'b01111; w[93][62] = 5'b00000; w[93][63] = 5'b10000; w[93][64] = 5'b01111; w[93][65] = 5'b01111; w[93][66] = 5'b01111; w[93][67] = 5'b00000; w[93][68] = 5'b01111; w[93][69] = 5'b01111; w[93][70] = 5'b01111; w[93][71] = 5'b01111; w[93][72] = 5'b00000; w[93][73] = 5'b01111; w[93][74] = 5'b01111; w[93][75] = 5'b01111; w[93][76] = 5'b00000; w[93][77] = 5'b10000; w[93][78] = 5'b01111; w[93][79] = 5'b01111; w[93][80] = 5'b01111; w[93][81] = 5'b00000; w[93][82] = 5'b01111; w[93][83] = 5'b01111; w[93][84] = 5'b01111; w[93][85] = 5'b01111; w[93][86] = 5'b00000; w[93][87] = 5'b01111; w[93][88] = 5'b01111; w[93][89] = 5'b01111; w[93][90] = 5'b00000; w[93][91] = 5'b00000; w[93][92] = 5'b01111; w[93][93] = 5'b00000; w[93][94] = 5'b01111; w[93][95] = 5'b01111; w[93][96] = 5'b01111; w[93][97] = 5'b01111; w[93][98] = 5'b01111; w[93][99] = 5'b01111; w[93][100] = 5'b00000; w[93][101] = 5'b01111; w[93][102] = 5'b01111; w[93][103] = 5'b01111; w[93][104] = 5'b00000; w[93][105] = 5'b00000; w[93][106] = 5'b00000; w[93][107] = 5'b01111; w[93][108] = 5'b01111; w[93][109] = 5'b00000; w[93][110] = 5'b01111; w[93][111] = 5'b01111; w[93][112] = 5'b01111; w[93][113] = 5'b01111; w[93][114] = 5'b00000; w[93][115] = 5'b01111; w[93][116] = 5'b01111; w[93][117] = 5'b01111; w[93][118] = 5'b00000; w[93][119] = 5'b00000; w[93][120] = 5'b01111; w[93][121] = 5'b01111; w[93][122] = 5'b01111; w[93][123] = 5'b00000; w[93][124] = 5'b01111; w[93][125] = 5'b01111; w[93][126] = 5'b01111; w[93][127] = 5'b01111; w[93][128] = 5'b00000; w[93][129] = 5'b01111; w[93][130] = 5'b01111; w[93][131] = 5'b01111; w[93][132] = 5'b10000; w[93][133] = 5'b00000; w[93][134] = 5'b01111; w[93][135] = 5'b01111; w[93][136] = 5'b01111; w[93][137] = 5'b00000; w[93][138] = 5'b01111; w[93][139] = 5'b01111; w[93][140] = 5'b01111; w[93][141] = 5'b01111; w[93][142] = 5'b00000; w[93][143] = 5'b01111; w[93][144] = 5'b01111; w[93][145] = 5'b01111; w[93][146] = 5'b10000; w[93][147] = 5'b00000; w[93][148] = 5'b01111; w[93][149] = 5'b01111; w[93][150] = 5'b01111; w[93][151] = 5'b00000; w[93][152] = 5'b01111; w[93][153] = 5'b01111; w[93][154] = 5'b01111; w[93][155] = 5'b01111; w[93][156] = 5'b01111; w[93][157] = 5'b01111; w[93][158] = 5'b01111; w[93][159] = 5'b10000; w[93][160] = 5'b10000; w[93][161] = 5'b10000; w[93][162] = 5'b00000; w[93][163] = 5'b01111; w[93][164] = 5'b01111; w[93][165] = 5'b01111; w[93][166] = 5'b01111; w[93][167] = 5'b01111; w[93][168] = 5'b01111; w[93][169] = 5'b01111; w[93][170] = 5'b01111; w[93][171] = 5'b01111; w[93][172] = 5'b01111; w[93][173] = 5'b10000; w[93][174] = 5'b10000; w[93][175] = 5'b10000; w[93][176] = 5'b00000; w[93][177] = 5'b01111; w[93][178] = 5'b01111; w[93][179] = 5'b01111; w[93][180] = 5'b01111; w[93][181] = 5'b01111; w[93][182] = 5'b01111; w[93][183] = 5'b01111; w[93][184] = 5'b01111; w[93][185] = 5'b01111; w[93][186] = 5'b01111; w[93][187] = 5'b01111; w[93][188] = 5'b01111; w[93][189] = 5'b01111; w[93][190] = 5'b01111; w[93][191] = 5'b01111; w[93][192] = 5'b01111; w[93][193] = 5'b01111; w[93][194] = 5'b01111; w[93][195] = 5'b01111; w[93][196] = 5'b01111; w[93][197] = 5'b01111; w[93][198] = 5'b01111; w[93][199] = 5'b01111; w[93][200] = 5'b01111; w[93][201] = 5'b01111; w[93][202] = 5'b01111; w[93][203] = 5'b01111; w[93][204] = 5'b01111; w[93][205] = 5'b01111; w[93][206] = 5'b01111; w[93][207] = 5'b01111; w[93][208] = 5'b01111; w[93][209] = 5'b01111; 
w[94][0] = 5'b01111; w[94][1] = 5'b01111; w[94][2] = 5'b01111; w[94][3] = 5'b01111; w[94][4] = 5'b01111; w[94][5] = 5'b01111; w[94][6] = 5'b01111; w[94][7] = 5'b01111; w[94][8] = 5'b01111; w[94][9] = 5'b01111; w[94][10] = 5'b01111; w[94][11] = 5'b01111; w[94][12] = 5'b01111; w[94][13] = 5'b01111; w[94][14] = 5'b01111; w[94][15] = 5'b01111; w[94][16] = 5'b01111; w[94][17] = 5'b01111; w[94][18] = 5'b01111; w[94][19] = 5'b01111; w[94][20] = 5'b01111; w[94][21] = 5'b01111; w[94][22] = 5'b01111; w[94][23] = 5'b01111; w[94][24] = 5'b01111; w[94][25] = 5'b01111; w[94][26] = 5'b01111; w[94][27] = 5'b01111; w[94][28] = 5'b01111; w[94][29] = 5'b01111; w[94][30] = 5'b00000; w[94][31] = 5'b01111; w[94][32] = 5'b00000; w[94][33] = 5'b10000; w[94][34] = 5'b10000; w[94][35] = 5'b10000; w[94][36] = 5'b10000; w[94][37] = 5'b00000; w[94][38] = 5'b01111; w[94][39] = 5'b00000; w[94][40] = 5'b01111; w[94][41] = 5'b01111; w[94][42] = 5'b01111; w[94][43] = 5'b01111; w[94][44] = 5'b00000; w[94][45] = 5'b00000; w[94][46] = 5'b00000; w[94][47] = 5'b10000; w[94][48] = 5'b10000; w[94][49] = 5'b10000; w[94][50] = 5'b10000; w[94][51] = 5'b00000; w[94][52] = 5'b00000; w[94][53] = 5'b00000; w[94][54] = 5'b01111; w[94][55] = 5'b01111; w[94][56] = 5'b01111; w[94][57] = 5'b01111; w[94][58] = 5'b00000; w[94][59] = 5'b01111; w[94][60] = 5'b01111; w[94][61] = 5'b01111; w[94][62] = 5'b00000; w[94][63] = 5'b10000; w[94][64] = 5'b01111; w[94][65] = 5'b01111; w[94][66] = 5'b01111; w[94][67] = 5'b00000; w[94][68] = 5'b01111; w[94][69] = 5'b01111; w[94][70] = 5'b01111; w[94][71] = 5'b01111; w[94][72] = 5'b00000; w[94][73] = 5'b01111; w[94][74] = 5'b01111; w[94][75] = 5'b01111; w[94][76] = 5'b00000; w[94][77] = 5'b10000; w[94][78] = 5'b01111; w[94][79] = 5'b01111; w[94][80] = 5'b01111; w[94][81] = 5'b00000; w[94][82] = 5'b01111; w[94][83] = 5'b01111; w[94][84] = 5'b01111; w[94][85] = 5'b01111; w[94][86] = 5'b00000; w[94][87] = 5'b01111; w[94][88] = 5'b01111; w[94][89] = 5'b01111; w[94][90] = 5'b00000; w[94][91] = 5'b00000; w[94][92] = 5'b01111; w[94][93] = 5'b01111; w[94][94] = 5'b00000; w[94][95] = 5'b01111; w[94][96] = 5'b01111; w[94][97] = 5'b01111; w[94][98] = 5'b01111; w[94][99] = 5'b01111; w[94][100] = 5'b00000; w[94][101] = 5'b01111; w[94][102] = 5'b01111; w[94][103] = 5'b01111; w[94][104] = 5'b00000; w[94][105] = 5'b00000; w[94][106] = 5'b00000; w[94][107] = 5'b01111; w[94][108] = 5'b01111; w[94][109] = 5'b00000; w[94][110] = 5'b01111; w[94][111] = 5'b01111; w[94][112] = 5'b01111; w[94][113] = 5'b01111; w[94][114] = 5'b00000; w[94][115] = 5'b01111; w[94][116] = 5'b01111; w[94][117] = 5'b01111; w[94][118] = 5'b00000; w[94][119] = 5'b00000; w[94][120] = 5'b01111; w[94][121] = 5'b01111; w[94][122] = 5'b01111; w[94][123] = 5'b00000; w[94][124] = 5'b01111; w[94][125] = 5'b01111; w[94][126] = 5'b01111; w[94][127] = 5'b01111; w[94][128] = 5'b00000; w[94][129] = 5'b01111; w[94][130] = 5'b01111; w[94][131] = 5'b01111; w[94][132] = 5'b10000; w[94][133] = 5'b00000; w[94][134] = 5'b01111; w[94][135] = 5'b01111; w[94][136] = 5'b01111; w[94][137] = 5'b00000; w[94][138] = 5'b01111; w[94][139] = 5'b01111; w[94][140] = 5'b01111; w[94][141] = 5'b01111; w[94][142] = 5'b00000; w[94][143] = 5'b01111; w[94][144] = 5'b01111; w[94][145] = 5'b01111; w[94][146] = 5'b10000; w[94][147] = 5'b00000; w[94][148] = 5'b01111; w[94][149] = 5'b01111; w[94][150] = 5'b01111; w[94][151] = 5'b00000; w[94][152] = 5'b01111; w[94][153] = 5'b01111; w[94][154] = 5'b01111; w[94][155] = 5'b01111; w[94][156] = 5'b01111; w[94][157] = 5'b01111; w[94][158] = 5'b01111; w[94][159] = 5'b10000; w[94][160] = 5'b10000; w[94][161] = 5'b10000; w[94][162] = 5'b00000; w[94][163] = 5'b01111; w[94][164] = 5'b01111; w[94][165] = 5'b01111; w[94][166] = 5'b01111; w[94][167] = 5'b01111; w[94][168] = 5'b01111; w[94][169] = 5'b01111; w[94][170] = 5'b01111; w[94][171] = 5'b01111; w[94][172] = 5'b01111; w[94][173] = 5'b10000; w[94][174] = 5'b10000; w[94][175] = 5'b10000; w[94][176] = 5'b00000; w[94][177] = 5'b01111; w[94][178] = 5'b01111; w[94][179] = 5'b01111; w[94][180] = 5'b01111; w[94][181] = 5'b01111; w[94][182] = 5'b01111; w[94][183] = 5'b01111; w[94][184] = 5'b01111; w[94][185] = 5'b01111; w[94][186] = 5'b01111; w[94][187] = 5'b01111; w[94][188] = 5'b01111; w[94][189] = 5'b01111; w[94][190] = 5'b01111; w[94][191] = 5'b01111; w[94][192] = 5'b01111; w[94][193] = 5'b01111; w[94][194] = 5'b01111; w[94][195] = 5'b01111; w[94][196] = 5'b01111; w[94][197] = 5'b01111; w[94][198] = 5'b01111; w[94][199] = 5'b01111; w[94][200] = 5'b01111; w[94][201] = 5'b01111; w[94][202] = 5'b01111; w[94][203] = 5'b01111; w[94][204] = 5'b01111; w[94][205] = 5'b01111; w[94][206] = 5'b01111; w[94][207] = 5'b01111; w[94][208] = 5'b01111; w[94][209] = 5'b01111; 
w[95][0] = 5'b01111; w[95][1] = 5'b01111; w[95][2] = 5'b01111; w[95][3] = 5'b01111; w[95][4] = 5'b01111; w[95][5] = 5'b01111; w[95][6] = 5'b01111; w[95][7] = 5'b01111; w[95][8] = 5'b01111; w[95][9] = 5'b01111; w[95][10] = 5'b01111; w[95][11] = 5'b01111; w[95][12] = 5'b01111; w[95][13] = 5'b01111; w[95][14] = 5'b01111; w[95][15] = 5'b01111; w[95][16] = 5'b01111; w[95][17] = 5'b01111; w[95][18] = 5'b01111; w[95][19] = 5'b01111; w[95][20] = 5'b01111; w[95][21] = 5'b01111; w[95][22] = 5'b01111; w[95][23] = 5'b01111; w[95][24] = 5'b01111; w[95][25] = 5'b01111; w[95][26] = 5'b01111; w[95][27] = 5'b01111; w[95][28] = 5'b01111; w[95][29] = 5'b01111; w[95][30] = 5'b01111; w[95][31] = 5'b00000; w[95][32] = 5'b10000; w[95][33] = 5'b10000; w[95][34] = 5'b10000; w[95][35] = 5'b10000; w[95][36] = 5'b10000; w[95][37] = 5'b10000; w[95][38] = 5'b00000; w[95][39] = 5'b01111; w[95][40] = 5'b01111; w[95][41] = 5'b01111; w[95][42] = 5'b01111; w[95][43] = 5'b01111; w[95][44] = 5'b01111; w[95][45] = 5'b10000; w[95][46] = 5'b10000; w[95][47] = 5'b10000; w[95][48] = 5'b10000; w[95][49] = 5'b10000; w[95][50] = 5'b10000; w[95][51] = 5'b10000; w[95][52] = 5'b10000; w[95][53] = 5'b01111; w[95][54] = 5'b01111; w[95][55] = 5'b01111; w[95][56] = 5'b01111; w[95][57] = 5'b01111; w[95][58] = 5'b01111; w[95][59] = 5'b00000; w[95][60] = 5'b00000; w[95][61] = 5'b01111; w[95][62] = 5'b10000; w[95][63] = 5'b00000; w[95][64] = 5'b01111; w[95][65] = 5'b00000; w[95][66] = 5'b00000; w[95][67] = 5'b01111; w[95][68] = 5'b01111; w[95][69] = 5'b01111; w[95][70] = 5'b01111; w[95][71] = 5'b01111; w[95][72] = 5'b01111; w[95][73] = 5'b00000; w[95][74] = 5'b01111; w[95][75] = 5'b01111; w[95][76] = 5'b10000; w[95][77] = 5'b00000; w[95][78] = 5'b01111; w[95][79] = 5'b01111; w[95][80] = 5'b00000; w[95][81] = 5'b01111; w[95][82] = 5'b01111; w[95][83] = 5'b01111; w[95][84] = 5'b01111; w[95][85] = 5'b01111; w[95][86] = 5'b01111; w[95][87] = 5'b00000; w[95][88] = 5'b01111; w[95][89] = 5'b01111; w[95][90] = 5'b10000; w[95][91] = 5'b10000; w[95][92] = 5'b01111; w[95][93] = 5'b01111; w[95][94] = 5'b01111; w[95][95] = 5'b00000; w[95][96] = 5'b01111; w[95][97] = 5'b01111; w[95][98] = 5'b01111; w[95][99] = 5'b01111; w[95][100] = 5'b01111; w[95][101] = 5'b00000; w[95][102] = 5'b01111; w[95][103] = 5'b01111; w[95][104] = 5'b10000; w[95][105] = 5'b10000; w[95][106] = 5'b01111; w[95][107] = 5'b00000; w[95][108] = 5'b00000; w[95][109] = 5'b01111; w[95][110] = 5'b01111; w[95][111] = 5'b01111; w[95][112] = 5'b01111; w[95][113] = 5'b01111; w[95][114] = 5'b01111; w[95][115] = 5'b00000; w[95][116] = 5'b01111; w[95][117] = 5'b01111; w[95][118] = 5'b10000; w[95][119] = 5'b10000; w[95][120] = 5'b00000; w[95][121] = 5'b00000; w[95][122] = 5'b00000; w[95][123] = 5'b01111; w[95][124] = 5'b01111; w[95][125] = 5'b01111; w[95][126] = 5'b01111; w[95][127] = 5'b01111; w[95][128] = 5'b01111; w[95][129] = 5'b00000; w[95][130] = 5'b01111; w[95][131] = 5'b01111; w[95][132] = 5'b00000; w[95][133] = 5'b10000; w[95][134] = 5'b01111; w[95][135] = 5'b01111; w[95][136] = 5'b00000; w[95][137] = 5'b01111; w[95][138] = 5'b01111; w[95][139] = 5'b01111; w[95][140] = 5'b01111; w[95][141] = 5'b01111; w[95][142] = 5'b01111; w[95][143] = 5'b00000; w[95][144] = 5'b00000; w[95][145] = 5'b01111; w[95][146] = 5'b00000; w[95][147] = 5'b10000; w[95][148] = 5'b01111; w[95][149] = 5'b00000; w[95][150] = 5'b00000; w[95][151] = 5'b01111; w[95][152] = 5'b01111; w[95][153] = 5'b01111; w[95][154] = 5'b01111; w[95][155] = 5'b01111; w[95][156] = 5'b01111; w[95][157] = 5'b00000; w[95][158] = 5'b00000; w[95][159] = 5'b00000; w[95][160] = 5'b10000; w[95][161] = 5'b10000; w[95][162] = 5'b10000; w[95][163] = 5'b00000; w[95][164] = 5'b00000; w[95][165] = 5'b01111; w[95][166] = 5'b01111; w[95][167] = 5'b01111; w[95][168] = 5'b01111; w[95][169] = 5'b01111; w[95][170] = 5'b01111; w[95][171] = 5'b01111; w[95][172] = 5'b00000; w[95][173] = 5'b00000; w[95][174] = 5'b10000; w[95][175] = 5'b10000; w[95][176] = 5'b10000; w[95][177] = 5'b00000; w[95][178] = 5'b01111; w[95][179] = 5'b01111; w[95][180] = 5'b01111; w[95][181] = 5'b01111; w[95][182] = 5'b01111; w[95][183] = 5'b01111; w[95][184] = 5'b01111; w[95][185] = 5'b01111; w[95][186] = 5'b01111; w[95][187] = 5'b01111; w[95][188] = 5'b01111; w[95][189] = 5'b01111; w[95][190] = 5'b01111; w[95][191] = 5'b01111; w[95][192] = 5'b01111; w[95][193] = 5'b01111; w[95][194] = 5'b01111; w[95][195] = 5'b01111; w[95][196] = 5'b01111; w[95][197] = 5'b01111; w[95][198] = 5'b01111; w[95][199] = 5'b01111; w[95][200] = 5'b01111; w[95][201] = 5'b01111; w[95][202] = 5'b01111; w[95][203] = 5'b01111; w[95][204] = 5'b01111; w[95][205] = 5'b01111; w[95][206] = 5'b01111; w[95][207] = 5'b01111; w[95][208] = 5'b01111; w[95][209] = 5'b01111; 
w[96][0] = 5'b01111; w[96][1] = 5'b01111; w[96][2] = 5'b01111; w[96][3] = 5'b01111; w[96][4] = 5'b01111; w[96][5] = 5'b01111; w[96][6] = 5'b01111; w[96][7] = 5'b01111; w[96][8] = 5'b01111; w[96][9] = 5'b01111; w[96][10] = 5'b01111; w[96][11] = 5'b01111; w[96][12] = 5'b01111; w[96][13] = 5'b01111; w[96][14] = 5'b01111; w[96][15] = 5'b01111; w[96][16] = 5'b01111; w[96][17] = 5'b01111; w[96][18] = 5'b01111; w[96][19] = 5'b01111; w[96][20] = 5'b01111; w[96][21] = 5'b01111; w[96][22] = 5'b01111; w[96][23] = 5'b01111; w[96][24] = 5'b01111; w[96][25] = 5'b01111; w[96][26] = 5'b01111; w[96][27] = 5'b01111; w[96][28] = 5'b01111; w[96][29] = 5'b01111; w[96][30] = 5'b01111; w[96][31] = 5'b00000; w[96][32] = 5'b10000; w[96][33] = 5'b10000; w[96][34] = 5'b10000; w[96][35] = 5'b10000; w[96][36] = 5'b10000; w[96][37] = 5'b10000; w[96][38] = 5'b00000; w[96][39] = 5'b01111; w[96][40] = 5'b01111; w[96][41] = 5'b01111; w[96][42] = 5'b01111; w[96][43] = 5'b01111; w[96][44] = 5'b01111; w[96][45] = 5'b10000; w[96][46] = 5'b10000; w[96][47] = 5'b10000; w[96][48] = 5'b10000; w[96][49] = 5'b10000; w[96][50] = 5'b10000; w[96][51] = 5'b10000; w[96][52] = 5'b10000; w[96][53] = 5'b01111; w[96][54] = 5'b01111; w[96][55] = 5'b01111; w[96][56] = 5'b01111; w[96][57] = 5'b01111; w[96][58] = 5'b01111; w[96][59] = 5'b00000; w[96][60] = 5'b00000; w[96][61] = 5'b01111; w[96][62] = 5'b10000; w[96][63] = 5'b00000; w[96][64] = 5'b01111; w[96][65] = 5'b00000; w[96][66] = 5'b00000; w[96][67] = 5'b01111; w[96][68] = 5'b01111; w[96][69] = 5'b01111; w[96][70] = 5'b01111; w[96][71] = 5'b01111; w[96][72] = 5'b01111; w[96][73] = 5'b00000; w[96][74] = 5'b01111; w[96][75] = 5'b01111; w[96][76] = 5'b10000; w[96][77] = 5'b00000; w[96][78] = 5'b01111; w[96][79] = 5'b01111; w[96][80] = 5'b00000; w[96][81] = 5'b01111; w[96][82] = 5'b01111; w[96][83] = 5'b01111; w[96][84] = 5'b01111; w[96][85] = 5'b01111; w[96][86] = 5'b01111; w[96][87] = 5'b00000; w[96][88] = 5'b01111; w[96][89] = 5'b01111; w[96][90] = 5'b10000; w[96][91] = 5'b10000; w[96][92] = 5'b01111; w[96][93] = 5'b01111; w[96][94] = 5'b01111; w[96][95] = 5'b01111; w[96][96] = 5'b00000; w[96][97] = 5'b01111; w[96][98] = 5'b01111; w[96][99] = 5'b01111; w[96][100] = 5'b01111; w[96][101] = 5'b00000; w[96][102] = 5'b01111; w[96][103] = 5'b01111; w[96][104] = 5'b10000; w[96][105] = 5'b10000; w[96][106] = 5'b01111; w[96][107] = 5'b00000; w[96][108] = 5'b00000; w[96][109] = 5'b01111; w[96][110] = 5'b01111; w[96][111] = 5'b01111; w[96][112] = 5'b01111; w[96][113] = 5'b01111; w[96][114] = 5'b01111; w[96][115] = 5'b00000; w[96][116] = 5'b01111; w[96][117] = 5'b01111; w[96][118] = 5'b10000; w[96][119] = 5'b10000; w[96][120] = 5'b00000; w[96][121] = 5'b00000; w[96][122] = 5'b00000; w[96][123] = 5'b01111; w[96][124] = 5'b01111; w[96][125] = 5'b01111; w[96][126] = 5'b01111; w[96][127] = 5'b01111; w[96][128] = 5'b01111; w[96][129] = 5'b00000; w[96][130] = 5'b01111; w[96][131] = 5'b01111; w[96][132] = 5'b00000; w[96][133] = 5'b10000; w[96][134] = 5'b01111; w[96][135] = 5'b01111; w[96][136] = 5'b00000; w[96][137] = 5'b01111; w[96][138] = 5'b01111; w[96][139] = 5'b01111; w[96][140] = 5'b01111; w[96][141] = 5'b01111; w[96][142] = 5'b01111; w[96][143] = 5'b00000; w[96][144] = 5'b00000; w[96][145] = 5'b01111; w[96][146] = 5'b00000; w[96][147] = 5'b10000; w[96][148] = 5'b01111; w[96][149] = 5'b00000; w[96][150] = 5'b00000; w[96][151] = 5'b01111; w[96][152] = 5'b01111; w[96][153] = 5'b01111; w[96][154] = 5'b01111; w[96][155] = 5'b01111; w[96][156] = 5'b01111; w[96][157] = 5'b00000; w[96][158] = 5'b00000; w[96][159] = 5'b00000; w[96][160] = 5'b10000; w[96][161] = 5'b10000; w[96][162] = 5'b10000; w[96][163] = 5'b00000; w[96][164] = 5'b00000; w[96][165] = 5'b01111; w[96][166] = 5'b01111; w[96][167] = 5'b01111; w[96][168] = 5'b01111; w[96][169] = 5'b01111; w[96][170] = 5'b01111; w[96][171] = 5'b01111; w[96][172] = 5'b00000; w[96][173] = 5'b00000; w[96][174] = 5'b10000; w[96][175] = 5'b10000; w[96][176] = 5'b10000; w[96][177] = 5'b00000; w[96][178] = 5'b01111; w[96][179] = 5'b01111; w[96][180] = 5'b01111; w[96][181] = 5'b01111; w[96][182] = 5'b01111; w[96][183] = 5'b01111; w[96][184] = 5'b01111; w[96][185] = 5'b01111; w[96][186] = 5'b01111; w[96][187] = 5'b01111; w[96][188] = 5'b01111; w[96][189] = 5'b01111; w[96][190] = 5'b01111; w[96][191] = 5'b01111; w[96][192] = 5'b01111; w[96][193] = 5'b01111; w[96][194] = 5'b01111; w[96][195] = 5'b01111; w[96][196] = 5'b01111; w[96][197] = 5'b01111; w[96][198] = 5'b01111; w[96][199] = 5'b01111; w[96][200] = 5'b01111; w[96][201] = 5'b01111; w[96][202] = 5'b01111; w[96][203] = 5'b01111; w[96][204] = 5'b01111; w[96][205] = 5'b01111; w[96][206] = 5'b01111; w[96][207] = 5'b01111; w[96][208] = 5'b01111; w[96][209] = 5'b01111; 
w[97][0] = 5'b01111; w[97][1] = 5'b01111; w[97][2] = 5'b01111; w[97][3] = 5'b01111; w[97][4] = 5'b01111; w[97][5] = 5'b01111; w[97][6] = 5'b01111; w[97][7] = 5'b01111; w[97][8] = 5'b01111; w[97][9] = 5'b01111; w[97][10] = 5'b01111; w[97][11] = 5'b01111; w[97][12] = 5'b01111; w[97][13] = 5'b01111; w[97][14] = 5'b01111; w[97][15] = 5'b01111; w[97][16] = 5'b01111; w[97][17] = 5'b01111; w[97][18] = 5'b01111; w[97][19] = 5'b01111; w[97][20] = 5'b01111; w[97][21] = 5'b01111; w[97][22] = 5'b01111; w[97][23] = 5'b01111; w[97][24] = 5'b01111; w[97][25] = 5'b01111; w[97][26] = 5'b01111; w[97][27] = 5'b01111; w[97][28] = 5'b01111; w[97][29] = 5'b01111; w[97][30] = 5'b01111; w[97][31] = 5'b00000; w[97][32] = 5'b10000; w[97][33] = 5'b10000; w[97][34] = 5'b10000; w[97][35] = 5'b10000; w[97][36] = 5'b10000; w[97][37] = 5'b10000; w[97][38] = 5'b00000; w[97][39] = 5'b01111; w[97][40] = 5'b01111; w[97][41] = 5'b01111; w[97][42] = 5'b01111; w[97][43] = 5'b01111; w[97][44] = 5'b01111; w[97][45] = 5'b10000; w[97][46] = 5'b10000; w[97][47] = 5'b10000; w[97][48] = 5'b10000; w[97][49] = 5'b10000; w[97][50] = 5'b10000; w[97][51] = 5'b10000; w[97][52] = 5'b10000; w[97][53] = 5'b01111; w[97][54] = 5'b01111; w[97][55] = 5'b01111; w[97][56] = 5'b01111; w[97][57] = 5'b01111; w[97][58] = 5'b01111; w[97][59] = 5'b00000; w[97][60] = 5'b00000; w[97][61] = 5'b01111; w[97][62] = 5'b10000; w[97][63] = 5'b00000; w[97][64] = 5'b01111; w[97][65] = 5'b00000; w[97][66] = 5'b00000; w[97][67] = 5'b01111; w[97][68] = 5'b01111; w[97][69] = 5'b01111; w[97][70] = 5'b01111; w[97][71] = 5'b01111; w[97][72] = 5'b01111; w[97][73] = 5'b00000; w[97][74] = 5'b01111; w[97][75] = 5'b01111; w[97][76] = 5'b10000; w[97][77] = 5'b00000; w[97][78] = 5'b01111; w[97][79] = 5'b01111; w[97][80] = 5'b00000; w[97][81] = 5'b01111; w[97][82] = 5'b01111; w[97][83] = 5'b01111; w[97][84] = 5'b01111; w[97][85] = 5'b01111; w[97][86] = 5'b01111; w[97][87] = 5'b00000; w[97][88] = 5'b01111; w[97][89] = 5'b01111; w[97][90] = 5'b10000; w[97][91] = 5'b10000; w[97][92] = 5'b01111; w[97][93] = 5'b01111; w[97][94] = 5'b01111; w[97][95] = 5'b01111; w[97][96] = 5'b01111; w[97][97] = 5'b00000; w[97][98] = 5'b01111; w[97][99] = 5'b01111; w[97][100] = 5'b01111; w[97][101] = 5'b00000; w[97][102] = 5'b01111; w[97][103] = 5'b01111; w[97][104] = 5'b10000; w[97][105] = 5'b10000; w[97][106] = 5'b01111; w[97][107] = 5'b00000; w[97][108] = 5'b00000; w[97][109] = 5'b01111; w[97][110] = 5'b01111; w[97][111] = 5'b01111; w[97][112] = 5'b01111; w[97][113] = 5'b01111; w[97][114] = 5'b01111; w[97][115] = 5'b00000; w[97][116] = 5'b01111; w[97][117] = 5'b01111; w[97][118] = 5'b10000; w[97][119] = 5'b10000; w[97][120] = 5'b00000; w[97][121] = 5'b00000; w[97][122] = 5'b00000; w[97][123] = 5'b01111; w[97][124] = 5'b01111; w[97][125] = 5'b01111; w[97][126] = 5'b01111; w[97][127] = 5'b01111; w[97][128] = 5'b01111; w[97][129] = 5'b00000; w[97][130] = 5'b01111; w[97][131] = 5'b01111; w[97][132] = 5'b00000; w[97][133] = 5'b10000; w[97][134] = 5'b01111; w[97][135] = 5'b01111; w[97][136] = 5'b00000; w[97][137] = 5'b01111; w[97][138] = 5'b01111; w[97][139] = 5'b01111; w[97][140] = 5'b01111; w[97][141] = 5'b01111; w[97][142] = 5'b01111; w[97][143] = 5'b00000; w[97][144] = 5'b00000; w[97][145] = 5'b01111; w[97][146] = 5'b00000; w[97][147] = 5'b10000; w[97][148] = 5'b01111; w[97][149] = 5'b00000; w[97][150] = 5'b00000; w[97][151] = 5'b01111; w[97][152] = 5'b01111; w[97][153] = 5'b01111; w[97][154] = 5'b01111; w[97][155] = 5'b01111; w[97][156] = 5'b01111; w[97][157] = 5'b00000; w[97][158] = 5'b00000; w[97][159] = 5'b00000; w[97][160] = 5'b10000; w[97][161] = 5'b10000; w[97][162] = 5'b10000; w[97][163] = 5'b00000; w[97][164] = 5'b00000; w[97][165] = 5'b01111; w[97][166] = 5'b01111; w[97][167] = 5'b01111; w[97][168] = 5'b01111; w[97][169] = 5'b01111; w[97][170] = 5'b01111; w[97][171] = 5'b01111; w[97][172] = 5'b00000; w[97][173] = 5'b00000; w[97][174] = 5'b10000; w[97][175] = 5'b10000; w[97][176] = 5'b10000; w[97][177] = 5'b00000; w[97][178] = 5'b01111; w[97][179] = 5'b01111; w[97][180] = 5'b01111; w[97][181] = 5'b01111; w[97][182] = 5'b01111; w[97][183] = 5'b01111; w[97][184] = 5'b01111; w[97][185] = 5'b01111; w[97][186] = 5'b01111; w[97][187] = 5'b01111; w[97][188] = 5'b01111; w[97][189] = 5'b01111; w[97][190] = 5'b01111; w[97][191] = 5'b01111; w[97][192] = 5'b01111; w[97][193] = 5'b01111; w[97][194] = 5'b01111; w[97][195] = 5'b01111; w[97][196] = 5'b01111; w[97][197] = 5'b01111; w[97][198] = 5'b01111; w[97][199] = 5'b01111; w[97][200] = 5'b01111; w[97][201] = 5'b01111; w[97][202] = 5'b01111; w[97][203] = 5'b01111; w[97][204] = 5'b01111; w[97][205] = 5'b01111; w[97][206] = 5'b01111; w[97][207] = 5'b01111; w[97][208] = 5'b01111; w[97][209] = 5'b01111; 
w[98][0] = 5'b01111; w[98][1] = 5'b01111; w[98][2] = 5'b01111; w[98][3] = 5'b01111; w[98][4] = 5'b01111; w[98][5] = 5'b01111; w[98][6] = 5'b01111; w[98][7] = 5'b01111; w[98][8] = 5'b01111; w[98][9] = 5'b01111; w[98][10] = 5'b01111; w[98][11] = 5'b01111; w[98][12] = 5'b01111; w[98][13] = 5'b01111; w[98][14] = 5'b01111; w[98][15] = 5'b01111; w[98][16] = 5'b01111; w[98][17] = 5'b01111; w[98][18] = 5'b01111; w[98][19] = 5'b01111; w[98][20] = 5'b01111; w[98][21] = 5'b01111; w[98][22] = 5'b01111; w[98][23] = 5'b01111; w[98][24] = 5'b01111; w[98][25] = 5'b01111; w[98][26] = 5'b01111; w[98][27] = 5'b01111; w[98][28] = 5'b01111; w[98][29] = 5'b01111; w[98][30] = 5'b01111; w[98][31] = 5'b00000; w[98][32] = 5'b10000; w[98][33] = 5'b10000; w[98][34] = 5'b10000; w[98][35] = 5'b10000; w[98][36] = 5'b10000; w[98][37] = 5'b10000; w[98][38] = 5'b00000; w[98][39] = 5'b01111; w[98][40] = 5'b01111; w[98][41] = 5'b01111; w[98][42] = 5'b01111; w[98][43] = 5'b01111; w[98][44] = 5'b01111; w[98][45] = 5'b10000; w[98][46] = 5'b10000; w[98][47] = 5'b10000; w[98][48] = 5'b10000; w[98][49] = 5'b10000; w[98][50] = 5'b10000; w[98][51] = 5'b10000; w[98][52] = 5'b10000; w[98][53] = 5'b01111; w[98][54] = 5'b01111; w[98][55] = 5'b01111; w[98][56] = 5'b01111; w[98][57] = 5'b01111; w[98][58] = 5'b01111; w[98][59] = 5'b00000; w[98][60] = 5'b00000; w[98][61] = 5'b01111; w[98][62] = 5'b10000; w[98][63] = 5'b00000; w[98][64] = 5'b01111; w[98][65] = 5'b00000; w[98][66] = 5'b00000; w[98][67] = 5'b01111; w[98][68] = 5'b01111; w[98][69] = 5'b01111; w[98][70] = 5'b01111; w[98][71] = 5'b01111; w[98][72] = 5'b01111; w[98][73] = 5'b00000; w[98][74] = 5'b01111; w[98][75] = 5'b01111; w[98][76] = 5'b10000; w[98][77] = 5'b00000; w[98][78] = 5'b01111; w[98][79] = 5'b01111; w[98][80] = 5'b00000; w[98][81] = 5'b01111; w[98][82] = 5'b01111; w[98][83] = 5'b01111; w[98][84] = 5'b01111; w[98][85] = 5'b01111; w[98][86] = 5'b01111; w[98][87] = 5'b00000; w[98][88] = 5'b01111; w[98][89] = 5'b01111; w[98][90] = 5'b10000; w[98][91] = 5'b10000; w[98][92] = 5'b01111; w[98][93] = 5'b01111; w[98][94] = 5'b01111; w[98][95] = 5'b01111; w[98][96] = 5'b01111; w[98][97] = 5'b01111; w[98][98] = 5'b00000; w[98][99] = 5'b01111; w[98][100] = 5'b01111; w[98][101] = 5'b00000; w[98][102] = 5'b01111; w[98][103] = 5'b01111; w[98][104] = 5'b10000; w[98][105] = 5'b10000; w[98][106] = 5'b01111; w[98][107] = 5'b00000; w[98][108] = 5'b00000; w[98][109] = 5'b01111; w[98][110] = 5'b01111; w[98][111] = 5'b01111; w[98][112] = 5'b01111; w[98][113] = 5'b01111; w[98][114] = 5'b01111; w[98][115] = 5'b00000; w[98][116] = 5'b01111; w[98][117] = 5'b01111; w[98][118] = 5'b10000; w[98][119] = 5'b10000; w[98][120] = 5'b00000; w[98][121] = 5'b00000; w[98][122] = 5'b00000; w[98][123] = 5'b01111; w[98][124] = 5'b01111; w[98][125] = 5'b01111; w[98][126] = 5'b01111; w[98][127] = 5'b01111; w[98][128] = 5'b01111; w[98][129] = 5'b00000; w[98][130] = 5'b01111; w[98][131] = 5'b01111; w[98][132] = 5'b00000; w[98][133] = 5'b10000; w[98][134] = 5'b01111; w[98][135] = 5'b01111; w[98][136] = 5'b00000; w[98][137] = 5'b01111; w[98][138] = 5'b01111; w[98][139] = 5'b01111; w[98][140] = 5'b01111; w[98][141] = 5'b01111; w[98][142] = 5'b01111; w[98][143] = 5'b00000; w[98][144] = 5'b00000; w[98][145] = 5'b01111; w[98][146] = 5'b00000; w[98][147] = 5'b10000; w[98][148] = 5'b01111; w[98][149] = 5'b00000; w[98][150] = 5'b00000; w[98][151] = 5'b01111; w[98][152] = 5'b01111; w[98][153] = 5'b01111; w[98][154] = 5'b01111; w[98][155] = 5'b01111; w[98][156] = 5'b01111; w[98][157] = 5'b00000; w[98][158] = 5'b00000; w[98][159] = 5'b00000; w[98][160] = 5'b10000; w[98][161] = 5'b10000; w[98][162] = 5'b10000; w[98][163] = 5'b00000; w[98][164] = 5'b00000; w[98][165] = 5'b01111; w[98][166] = 5'b01111; w[98][167] = 5'b01111; w[98][168] = 5'b01111; w[98][169] = 5'b01111; w[98][170] = 5'b01111; w[98][171] = 5'b01111; w[98][172] = 5'b00000; w[98][173] = 5'b00000; w[98][174] = 5'b10000; w[98][175] = 5'b10000; w[98][176] = 5'b10000; w[98][177] = 5'b00000; w[98][178] = 5'b01111; w[98][179] = 5'b01111; w[98][180] = 5'b01111; w[98][181] = 5'b01111; w[98][182] = 5'b01111; w[98][183] = 5'b01111; w[98][184] = 5'b01111; w[98][185] = 5'b01111; w[98][186] = 5'b01111; w[98][187] = 5'b01111; w[98][188] = 5'b01111; w[98][189] = 5'b01111; w[98][190] = 5'b01111; w[98][191] = 5'b01111; w[98][192] = 5'b01111; w[98][193] = 5'b01111; w[98][194] = 5'b01111; w[98][195] = 5'b01111; w[98][196] = 5'b01111; w[98][197] = 5'b01111; w[98][198] = 5'b01111; w[98][199] = 5'b01111; w[98][200] = 5'b01111; w[98][201] = 5'b01111; w[98][202] = 5'b01111; w[98][203] = 5'b01111; w[98][204] = 5'b01111; w[98][205] = 5'b01111; w[98][206] = 5'b01111; w[98][207] = 5'b01111; w[98][208] = 5'b01111; w[98][209] = 5'b01111; 
w[99][0] = 5'b01111; w[99][1] = 5'b01111; w[99][2] = 5'b01111; w[99][3] = 5'b01111; w[99][4] = 5'b01111; w[99][5] = 5'b01111; w[99][6] = 5'b01111; w[99][7] = 5'b01111; w[99][8] = 5'b01111; w[99][9] = 5'b01111; w[99][10] = 5'b01111; w[99][11] = 5'b01111; w[99][12] = 5'b01111; w[99][13] = 5'b01111; w[99][14] = 5'b01111; w[99][15] = 5'b01111; w[99][16] = 5'b01111; w[99][17] = 5'b01111; w[99][18] = 5'b01111; w[99][19] = 5'b01111; w[99][20] = 5'b01111; w[99][21] = 5'b01111; w[99][22] = 5'b01111; w[99][23] = 5'b01111; w[99][24] = 5'b01111; w[99][25] = 5'b01111; w[99][26] = 5'b01111; w[99][27] = 5'b01111; w[99][28] = 5'b01111; w[99][29] = 5'b01111; w[99][30] = 5'b01111; w[99][31] = 5'b00000; w[99][32] = 5'b10000; w[99][33] = 5'b10000; w[99][34] = 5'b10000; w[99][35] = 5'b10000; w[99][36] = 5'b10000; w[99][37] = 5'b10000; w[99][38] = 5'b00000; w[99][39] = 5'b01111; w[99][40] = 5'b01111; w[99][41] = 5'b01111; w[99][42] = 5'b01111; w[99][43] = 5'b01111; w[99][44] = 5'b01111; w[99][45] = 5'b10000; w[99][46] = 5'b10000; w[99][47] = 5'b10000; w[99][48] = 5'b10000; w[99][49] = 5'b10000; w[99][50] = 5'b10000; w[99][51] = 5'b10000; w[99][52] = 5'b10000; w[99][53] = 5'b01111; w[99][54] = 5'b01111; w[99][55] = 5'b01111; w[99][56] = 5'b01111; w[99][57] = 5'b01111; w[99][58] = 5'b01111; w[99][59] = 5'b00000; w[99][60] = 5'b00000; w[99][61] = 5'b01111; w[99][62] = 5'b10000; w[99][63] = 5'b00000; w[99][64] = 5'b01111; w[99][65] = 5'b00000; w[99][66] = 5'b00000; w[99][67] = 5'b01111; w[99][68] = 5'b01111; w[99][69] = 5'b01111; w[99][70] = 5'b01111; w[99][71] = 5'b01111; w[99][72] = 5'b01111; w[99][73] = 5'b00000; w[99][74] = 5'b01111; w[99][75] = 5'b01111; w[99][76] = 5'b10000; w[99][77] = 5'b00000; w[99][78] = 5'b01111; w[99][79] = 5'b01111; w[99][80] = 5'b00000; w[99][81] = 5'b01111; w[99][82] = 5'b01111; w[99][83] = 5'b01111; w[99][84] = 5'b01111; w[99][85] = 5'b01111; w[99][86] = 5'b01111; w[99][87] = 5'b00000; w[99][88] = 5'b01111; w[99][89] = 5'b01111; w[99][90] = 5'b10000; w[99][91] = 5'b10000; w[99][92] = 5'b01111; w[99][93] = 5'b01111; w[99][94] = 5'b01111; w[99][95] = 5'b01111; w[99][96] = 5'b01111; w[99][97] = 5'b01111; w[99][98] = 5'b01111; w[99][99] = 5'b00000; w[99][100] = 5'b01111; w[99][101] = 5'b00000; w[99][102] = 5'b01111; w[99][103] = 5'b01111; w[99][104] = 5'b10000; w[99][105] = 5'b10000; w[99][106] = 5'b01111; w[99][107] = 5'b00000; w[99][108] = 5'b00000; w[99][109] = 5'b01111; w[99][110] = 5'b01111; w[99][111] = 5'b01111; w[99][112] = 5'b01111; w[99][113] = 5'b01111; w[99][114] = 5'b01111; w[99][115] = 5'b00000; w[99][116] = 5'b01111; w[99][117] = 5'b01111; w[99][118] = 5'b10000; w[99][119] = 5'b10000; w[99][120] = 5'b00000; w[99][121] = 5'b00000; w[99][122] = 5'b00000; w[99][123] = 5'b01111; w[99][124] = 5'b01111; w[99][125] = 5'b01111; w[99][126] = 5'b01111; w[99][127] = 5'b01111; w[99][128] = 5'b01111; w[99][129] = 5'b00000; w[99][130] = 5'b01111; w[99][131] = 5'b01111; w[99][132] = 5'b00000; w[99][133] = 5'b10000; w[99][134] = 5'b01111; w[99][135] = 5'b01111; w[99][136] = 5'b00000; w[99][137] = 5'b01111; w[99][138] = 5'b01111; w[99][139] = 5'b01111; w[99][140] = 5'b01111; w[99][141] = 5'b01111; w[99][142] = 5'b01111; w[99][143] = 5'b00000; w[99][144] = 5'b00000; w[99][145] = 5'b01111; w[99][146] = 5'b00000; w[99][147] = 5'b10000; w[99][148] = 5'b01111; w[99][149] = 5'b00000; w[99][150] = 5'b00000; w[99][151] = 5'b01111; w[99][152] = 5'b01111; w[99][153] = 5'b01111; w[99][154] = 5'b01111; w[99][155] = 5'b01111; w[99][156] = 5'b01111; w[99][157] = 5'b00000; w[99][158] = 5'b00000; w[99][159] = 5'b00000; w[99][160] = 5'b10000; w[99][161] = 5'b10000; w[99][162] = 5'b10000; w[99][163] = 5'b00000; w[99][164] = 5'b00000; w[99][165] = 5'b01111; w[99][166] = 5'b01111; w[99][167] = 5'b01111; w[99][168] = 5'b01111; w[99][169] = 5'b01111; w[99][170] = 5'b01111; w[99][171] = 5'b01111; w[99][172] = 5'b00000; w[99][173] = 5'b00000; w[99][174] = 5'b10000; w[99][175] = 5'b10000; w[99][176] = 5'b10000; w[99][177] = 5'b00000; w[99][178] = 5'b01111; w[99][179] = 5'b01111; w[99][180] = 5'b01111; w[99][181] = 5'b01111; w[99][182] = 5'b01111; w[99][183] = 5'b01111; w[99][184] = 5'b01111; w[99][185] = 5'b01111; w[99][186] = 5'b01111; w[99][187] = 5'b01111; w[99][188] = 5'b01111; w[99][189] = 5'b01111; w[99][190] = 5'b01111; w[99][191] = 5'b01111; w[99][192] = 5'b01111; w[99][193] = 5'b01111; w[99][194] = 5'b01111; w[99][195] = 5'b01111; w[99][196] = 5'b01111; w[99][197] = 5'b01111; w[99][198] = 5'b01111; w[99][199] = 5'b01111; w[99][200] = 5'b01111; w[99][201] = 5'b01111; w[99][202] = 5'b01111; w[99][203] = 5'b01111; w[99][204] = 5'b01111; w[99][205] = 5'b01111; w[99][206] = 5'b01111; w[99][207] = 5'b01111; w[99][208] = 5'b01111; w[99][209] = 5'b01111; 
w[100][0] = 5'b01111; w[100][1] = 5'b01111; w[100][2] = 5'b01111; w[100][3] = 5'b01111; w[100][4] = 5'b01111; w[100][5] = 5'b01111; w[100][6] = 5'b01111; w[100][7] = 5'b01111; w[100][8] = 5'b01111; w[100][9] = 5'b01111; w[100][10] = 5'b01111; w[100][11] = 5'b01111; w[100][12] = 5'b01111; w[100][13] = 5'b01111; w[100][14] = 5'b01111; w[100][15] = 5'b01111; w[100][16] = 5'b01111; w[100][17] = 5'b01111; w[100][18] = 5'b01111; w[100][19] = 5'b01111; w[100][20] = 5'b01111; w[100][21] = 5'b01111; w[100][22] = 5'b01111; w[100][23] = 5'b01111; w[100][24] = 5'b01111; w[100][25] = 5'b01111; w[100][26] = 5'b01111; w[100][27] = 5'b01111; w[100][28] = 5'b01111; w[100][29] = 5'b01111; w[100][30] = 5'b00000; w[100][31] = 5'b10000; w[100][32] = 5'b00000; w[100][33] = 5'b10000; w[100][34] = 5'b00000; w[100][35] = 5'b00000; w[100][36] = 5'b00000; w[100][37] = 5'b00000; w[100][38] = 5'b10000; w[100][39] = 5'b00000; w[100][40] = 5'b01111; w[100][41] = 5'b01111; w[100][42] = 5'b01111; w[100][43] = 5'b01111; w[100][44] = 5'b00000; w[100][45] = 5'b00000; w[100][46] = 5'b00000; w[100][47] = 5'b10000; w[100][48] = 5'b00000; w[100][49] = 5'b00000; w[100][50] = 5'b00000; w[100][51] = 5'b00000; w[100][52] = 5'b00000; w[100][53] = 5'b00000; w[100][54] = 5'b01111; w[100][55] = 5'b01111; w[100][56] = 5'b01111; w[100][57] = 5'b01111; w[100][58] = 5'b01111; w[100][59] = 5'b01111; w[100][60] = 5'b01111; w[100][61] = 5'b00000; w[100][62] = 5'b10000; w[100][63] = 5'b10000; w[100][64] = 5'b01111; w[100][65] = 5'b01111; w[100][66] = 5'b01111; w[100][67] = 5'b01111; w[100][68] = 5'b01111; w[100][69] = 5'b01111; w[100][70] = 5'b01111; w[100][71] = 5'b01111; w[100][72] = 5'b01111; w[100][73] = 5'b01111; w[100][74] = 5'b00000; w[100][75] = 5'b00000; w[100][76] = 5'b10000; w[100][77] = 5'b10000; w[100][78] = 5'b01111; w[100][79] = 5'b00000; w[100][80] = 5'b01111; w[100][81] = 5'b01111; w[100][82] = 5'b01111; w[100][83] = 5'b01111; w[100][84] = 5'b01111; w[100][85] = 5'b01111; w[100][86] = 5'b01111; w[100][87] = 5'b01111; w[100][88] = 5'b00000; w[100][89] = 5'b00000; w[100][90] = 5'b10000; w[100][91] = 5'b10000; w[100][92] = 5'b01111; w[100][93] = 5'b00000; w[100][94] = 5'b00000; w[100][95] = 5'b01111; w[100][96] = 5'b01111; w[100][97] = 5'b01111; w[100][98] = 5'b01111; w[100][99] = 5'b01111; w[100][100] = 5'b00000; w[100][101] = 5'b01111; w[100][102] = 5'b00000; w[100][103] = 5'b01111; w[100][104] = 5'b10000; w[100][105] = 5'b10000; w[100][106] = 5'b01111; w[100][107] = 5'b01111; w[100][108] = 5'b01111; w[100][109] = 5'b01111; w[100][110] = 5'b01111; w[100][111] = 5'b01111; w[100][112] = 5'b01111; w[100][113] = 5'b01111; w[100][114] = 5'b01111; w[100][115] = 5'b01111; w[100][116] = 5'b00000; w[100][117] = 5'b01111; w[100][118] = 5'b10000; w[100][119] = 5'b10000; w[100][120] = 5'b01111; w[100][121] = 5'b01111; w[100][122] = 5'b01111; w[100][123] = 5'b01111; w[100][124] = 5'b01111; w[100][125] = 5'b01111; w[100][126] = 5'b01111; w[100][127] = 5'b01111; w[100][128] = 5'b01111; w[100][129] = 5'b01111; w[100][130] = 5'b00000; w[100][131] = 5'b01111; w[100][132] = 5'b10000; w[100][133] = 5'b10000; w[100][134] = 5'b00000; w[100][135] = 5'b00000; w[100][136] = 5'b01111; w[100][137] = 5'b01111; w[100][138] = 5'b01111; w[100][139] = 5'b01111; w[100][140] = 5'b01111; w[100][141] = 5'b01111; w[100][142] = 5'b01111; w[100][143] = 5'b01111; w[100][144] = 5'b01111; w[100][145] = 5'b01111; w[100][146] = 5'b10000; w[100][147] = 5'b10000; w[100][148] = 5'b00000; w[100][149] = 5'b01111; w[100][150] = 5'b01111; w[100][151] = 5'b01111; w[100][152] = 5'b01111; w[100][153] = 5'b01111; w[100][154] = 5'b01111; w[100][155] = 5'b01111; w[100][156] = 5'b01111; w[100][157] = 5'b01111; w[100][158] = 5'b01111; w[100][159] = 5'b01111; w[100][160] = 5'b00000; w[100][161] = 5'b00000; w[100][162] = 5'b00000; w[100][163] = 5'b01111; w[100][164] = 5'b01111; w[100][165] = 5'b01111; w[100][166] = 5'b01111; w[100][167] = 5'b01111; w[100][168] = 5'b01111; w[100][169] = 5'b01111; w[100][170] = 5'b01111; w[100][171] = 5'b00000; w[100][172] = 5'b01111; w[100][173] = 5'b01111; w[100][174] = 5'b00000; w[100][175] = 5'b00000; w[100][176] = 5'b00000; w[100][177] = 5'b01111; w[100][178] = 5'b00000; w[100][179] = 5'b01111; w[100][180] = 5'b01111; w[100][181] = 5'b01111; w[100][182] = 5'b01111; w[100][183] = 5'b01111; w[100][184] = 5'b01111; w[100][185] = 5'b01111; w[100][186] = 5'b01111; w[100][187] = 5'b01111; w[100][188] = 5'b01111; w[100][189] = 5'b01111; w[100][190] = 5'b01111; w[100][191] = 5'b01111; w[100][192] = 5'b01111; w[100][193] = 5'b01111; w[100][194] = 5'b01111; w[100][195] = 5'b01111; w[100][196] = 5'b01111; w[100][197] = 5'b01111; w[100][198] = 5'b01111; w[100][199] = 5'b01111; w[100][200] = 5'b01111; w[100][201] = 5'b01111; w[100][202] = 5'b01111; w[100][203] = 5'b01111; w[100][204] = 5'b01111; w[100][205] = 5'b01111; w[100][206] = 5'b01111; w[100][207] = 5'b01111; w[100][208] = 5'b01111; w[100][209] = 5'b01111; 
w[101][0] = 5'b00000; w[101][1] = 5'b00000; w[101][2] = 5'b00000; w[101][3] = 5'b00000; w[101][4] = 5'b00000; w[101][5] = 5'b00000; w[101][6] = 5'b00000; w[101][7] = 5'b00000; w[101][8] = 5'b00000; w[101][9] = 5'b00000; w[101][10] = 5'b00000; w[101][11] = 5'b00000; w[101][12] = 5'b00000; w[101][13] = 5'b00000; w[101][14] = 5'b00000; w[101][15] = 5'b00000; w[101][16] = 5'b00000; w[101][17] = 5'b00000; w[101][18] = 5'b00000; w[101][19] = 5'b00000; w[101][20] = 5'b00000; w[101][21] = 5'b00000; w[101][22] = 5'b00000; w[101][23] = 5'b00000; w[101][24] = 5'b00000; w[101][25] = 5'b00000; w[101][26] = 5'b00000; w[101][27] = 5'b00000; w[101][28] = 5'b00000; w[101][29] = 5'b00000; w[101][30] = 5'b10000; w[101][31] = 5'b00000; w[101][32] = 5'b01111; w[101][33] = 5'b00000; w[101][34] = 5'b10000; w[101][35] = 5'b10000; w[101][36] = 5'b10000; w[101][37] = 5'b01111; w[101][38] = 5'b00000; w[101][39] = 5'b10000; w[101][40] = 5'b00000; w[101][41] = 5'b00000; w[101][42] = 5'b00000; w[101][43] = 5'b00000; w[101][44] = 5'b10000; w[101][45] = 5'b01111; w[101][46] = 5'b01111; w[101][47] = 5'b00000; w[101][48] = 5'b10000; w[101][49] = 5'b10000; w[101][50] = 5'b10000; w[101][51] = 5'b01111; w[101][52] = 5'b01111; w[101][53] = 5'b10000; w[101][54] = 5'b00000; w[101][55] = 5'b00000; w[101][56] = 5'b00000; w[101][57] = 5'b00000; w[101][58] = 5'b01111; w[101][59] = 5'b01111; w[101][60] = 5'b01111; w[101][61] = 5'b01111; w[101][62] = 5'b10000; w[101][63] = 5'b10000; w[101][64] = 5'b00000; w[101][65] = 5'b01111; w[101][66] = 5'b01111; w[101][67] = 5'b01111; w[101][68] = 5'b00000; w[101][69] = 5'b00000; w[101][70] = 5'b00000; w[101][71] = 5'b00000; w[101][72] = 5'b01111; w[101][73] = 5'b01111; w[101][74] = 5'b01111; w[101][75] = 5'b01111; w[101][76] = 5'b10000; w[101][77] = 5'b10000; w[101][78] = 5'b00000; w[101][79] = 5'b01111; w[101][80] = 5'b01111; w[101][81] = 5'b01111; w[101][82] = 5'b00000; w[101][83] = 5'b00000; w[101][84] = 5'b00000; w[101][85] = 5'b00000; w[101][86] = 5'b01111; w[101][87] = 5'b01111; w[101][88] = 5'b01111; w[101][89] = 5'b01111; w[101][90] = 5'b10000; w[101][91] = 5'b10000; w[101][92] = 5'b00000; w[101][93] = 5'b01111; w[101][94] = 5'b01111; w[101][95] = 5'b00000; w[101][96] = 5'b00000; w[101][97] = 5'b00000; w[101][98] = 5'b00000; w[101][99] = 5'b00000; w[101][100] = 5'b01111; w[101][101] = 5'b00000; w[101][102] = 5'b01111; w[101][103] = 5'b00000; w[101][104] = 5'b10000; w[101][105] = 5'b10000; w[101][106] = 5'b01111; w[101][107] = 5'b01111; w[101][108] = 5'b01111; w[101][109] = 5'b01111; w[101][110] = 5'b00000; w[101][111] = 5'b00000; w[101][112] = 5'b00000; w[101][113] = 5'b00000; w[101][114] = 5'b01111; w[101][115] = 5'b01111; w[101][116] = 5'b01111; w[101][117] = 5'b00000; w[101][118] = 5'b10000; w[101][119] = 5'b10000; w[101][120] = 5'b01111; w[101][121] = 5'b01111; w[101][122] = 5'b01111; w[101][123] = 5'b01111; w[101][124] = 5'b00000; w[101][125] = 5'b00000; w[101][126] = 5'b00000; w[101][127] = 5'b00000; w[101][128] = 5'b01111; w[101][129] = 5'b01111; w[101][130] = 5'b01111; w[101][131] = 5'b00000; w[101][132] = 5'b10000; w[101][133] = 5'b10000; w[101][134] = 5'b01111; w[101][135] = 5'b01111; w[101][136] = 5'b01111; w[101][137] = 5'b01111; w[101][138] = 5'b00000; w[101][139] = 5'b00000; w[101][140] = 5'b00000; w[101][141] = 5'b00000; w[101][142] = 5'b01111; w[101][143] = 5'b01111; w[101][144] = 5'b01111; w[101][145] = 5'b00000; w[101][146] = 5'b10000; w[101][147] = 5'b10000; w[101][148] = 5'b01111; w[101][149] = 5'b01111; w[101][150] = 5'b01111; w[101][151] = 5'b01111; w[101][152] = 5'b00000; w[101][153] = 5'b00000; w[101][154] = 5'b00000; w[101][155] = 5'b00000; w[101][156] = 5'b00000; w[101][157] = 5'b01111; w[101][158] = 5'b01111; w[101][159] = 5'b00000; w[101][160] = 5'b10000; w[101][161] = 5'b10000; w[101][162] = 5'b01111; w[101][163] = 5'b01111; w[101][164] = 5'b01111; w[101][165] = 5'b00000; w[101][166] = 5'b00000; w[101][167] = 5'b00000; w[101][168] = 5'b00000; w[101][169] = 5'b00000; w[101][170] = 5'b00000; w[101][171] = 5'b01111; w[101][172] = 5'b01111; w[101][173] = 5'b00000; w[101][174] = 5'b10000; w[101][175] = 5'b10000; w[101][176] = 5'b01111; w[101][177] = 5'b01111; w[101][178] = 5'b01111; w[101][179] = 5'b00000; w[101][180] = 5'b00000; w[101][181] = 5'b00000; w[101][182] = 5'b00000; w[101][183] = 5'b00000; w[101][184] = 5'b00000; w[101][185] = 5'b00000; w[101][186] = 5'b00000; w[101][187] = 5'b00000; w[101][188] = 5'b00000; w[101][189] = 5'b00000; w[101][190] = 5'b00000; w[101][191] = 5'b00000; w[101][192] = 5'b00000; w[101][193] = 5'b00000; w[101][194] = 5'b00000; w[101][195] = 5'b00000; w[101][196] = 5'b00000; w[101][197] = 5'b00000; w[101][198] = 5'b00000; w[101][199] = 5'b00000; w[101][200] = 5'b00000; w[101][201] = 5'b00000; w[101][202] = 5'b00000; w[101][203] = 5'b00000; w[101][204] = 5'b00000; w[101][205] = 5'b00000; w[101][206] = 5'b00000; w[101][207] = 5'b00000; w[101][208] = 5'b00000; w[101][209] = 5'b00000; 
w[102][0] = 5'b01111; w[102][1] = 5'b01111; w[102][2] = 5'b01111; w[102][3] = 5'b01111; w[102][4] = 5'b01111; w[102][5] = 5'b01111; w[102][6] = 5'b01111; w[102][7] = 5'b01111; w[102][8] = 5'b01111; w[102][9] = 5'b01111; w[102][10] = 5'b01111; w[102][11] = 5'b01111; w[102][12] = 5'b01111; w[102][13] = 5'b01111; w[102][14] = 5'b01111; w[102][15] = 5'b01111; w[102][16] = 5'b01111; w[102][17] = 5'b01111; w[102][18] = 5'b01111; w[102][19] = 5'b01111; w[102][20] = 5'b01111; w[102][21] = 5'b01111; w[102][22] = 5'b01111; w[102][23] = 5'b01111; w[102][24] = 5'b01111; w[102][25] = 5'b01111; w[102][26] = 5'b01111; w[102][27] = 5'b01111; w[102][28] = 5'b01111; w[102][29] = 5'b01111; w[102][30] = 5'b00000; w[102][31] = 5'b01111; w[102][32] = 5'b00000; w[102][33] = 5'b10000; w[102][34] = 5'b10000; w[102][35] = 5'b10000; w[102][36] = 5'b10000; w[102][37] = 5'b00000; w[102][38] = 5'b01111; w[102][39] = 5'b00000; w[102][40] = 5'b01111; w[102][41] = 5'b01111; w[102][42] = 5'b01111; w[102][43] = 5'b01111; w[102][44] = 5'b00000; w[102][45] = 5'b00000; w[102][46] = 5'b00000; w[102][47] = 5'b10000; w[102][48] = 5'b10000; w[102][49] = 5'b10000; w[102][50] = 5'b10000; w[102][51] = 5'b00000; w[102][52] = 5'b00000; w[102][53] = 5'b00000; w[102][54] = 5'b01111; w[102][55] = 5'b01111; w[102][56] = 5'b01111; w[102][57] = 5'b01111; w[102][58] = 5'b00000; w[102][59] = 5'b01111; w[102][60] = 5'b01111; w[102][61] = 5'b01111; w[102][62] = 5'b00000; w[102][63] = 5'b10000; w[102][64] = 5'b01111; w[102][65] = 5'b01111; w[102][66] = 5'b01111; w[102][67] = 5'b00000; w[102][68] = 5'b01111; w[102][69] = 5'b01111; w[102][70] = 5'b01111; w[102][71] = 5'b01111; w[102][72] = 5'b00000; w[102][73] = 5'b01111; w[102][74] = 5'b01111; w[102][75] = 5'b01111; w[102][76] = 5'b00000; w[102][77] = 5'b10000; w[102][78] = 5'b01111; w[102][79] = 5'b01111; w[102][80] = 5'b01111; w[102][81] = 5'b00000; w[102][82] = 5'b01111; w[102][83] = 5'b01111; w[102][84] = 5'b01111; w[102][85] = 5'b01111; w[102][86] = 5'b00000; w[102][87] = 5'b01111; w[102][88] = 5'b01111; w[102][89] = 5'b01111; w[102][90] = 5'b00000; w[102][91] = 5'b00000; w[102][92] = 5'b01111; w[102][93] = 5'b01111; w[102][94] = 5'b01111; w[102][95] = 5'b01111; w[102][96] = 5'b01111; w[102][97] = 5'b01111; w[102][98] = 5'b01111; w[102][99] = 5'b01111; w[102][100] = 5'b00000; w[102][101] = 5'b01111; w[102][102] = 5'b00000; w[102][103] = 5'b01111; w[102][104] = 5'b00000; w[102][105] = 5'b00000; w[102][106] = 5'b00000; w[102][107] = 5'b01111; w[102][108] = 5'b01111; w[102][109] = 5'b00000; w[102][110] = 5'b01111; w[102][111] = 5'b01111; w[102][112] = 5'b01111; w[102][113] = 5'b01111; w[102][114] = 5'b00000; w[102][115] = 5'b01111; w[102][116] = 5'b01111; w[102][117] = 5'b01111; w[102][118] = 5'b00000; w[102][119] = 5'b00000; w[102][120] = 5'b01111; w[102][121] = 5'b01111; w[102][122] = 5'b01111; w[102][123] = 5'b00000; w[102][124] = 5'b01111; w[102][125] = 5'b01111; w[102][126] = 5'b01111; w[102][127] = 5'b01111; w[102][128] = 5'b00000; w[102][129] = 5'b01111; w[102][130] = 5'b01111; w[102][131] = 5'b01111; w[102][132] = 5'b10000; w[102][133] = 5'b00000; w[102][134] = 5'b01111; w[102][135] = 5'b01111; w[102][136] = 5'b01111; w[102][137] = 5'b00000; w[102][138] = 5'b01111; w[102][139] = 5'b01111; w[102][140] = 5'b01111; w[102][141] = 5'b01111; w[102][142] = 5'b00000; w[102][143] = 5'b01111; w[102][144] = 5'b01111; w[102][145] = 5'b01111; w[102][146] = 5'b10000; w[102][147] = 5'b00000; w[102][148] = 5'b01111; w[102][149] = 5'b01111; w[102][150] = 5'b01111; w[102][151] = 5'b00000; w[102][152] = 5'b01111; w[102][153] = 5'b01111; w[102][154] = 5'b01111; w[102][155] = 5'b01111; w[102][156] = 5'b01111; w[102][157] = 5'b01111; w[102][158] = 5'b01111; w[102][159] = 5'b10000; w[102][160] = 5'b10000; w[102][161] = 5'b10000; w[102][162] = 5'b00000; w[102][163] = 5'b01111; w[102][164] = 5'b01111; w[102][165] = 5'b01111; w[102][166] = 5'b01111; w[102][167] = 5'b01111; w[102][168] = 5'b01111; w[102][169] = 5'b01111; w[102][170] = 5'b01111; w[102][171] = 5'b01111; w[102][172] = 5'b01111; w[102][173] = 5'b10000; w[102][174] = 5'b10000; w[102][175] = 5'b10000; w[102][176] = 5'b00000; w[102][177] = 5'b01111; w[102][178] = 5'b01111; w[102][179] = 5'b01111; w[102][180] = 5'b01111; w[102][181] = 5'b01111; w[102][182] = 5'b01111; w[102][183] = 5'b01111; w[102][184] = 5'b01111; w[102][185] = 5'b01111; w[102][186] = 5'b01111; w[102][187] = 5'b01111; w[102][188] = 5'b01111; w[102][189] = 5'b01111; w[102][190] = 5'b01111; w[102][191] = 5'b01111; w[102][192] = 5'b01111; w[102][193] = 5'b01111; w[102][194] = 5'b01111; w[102][195] = 5'b01111; w[102][196] = 5'b01111; w[102][197] = 5'b01111; w[102][198] = 5'b01111; w[102][199] = 5'b01111; w[102][200] = 5'b01111; w[102][201] = 5'b01111; w[102][202] = 5'b01111; w[102][203] = 5'b01111; w[102][204] = 5'b01111; w[102][205] = 5'b01111; w[102][206] = 5'b01111; w[102][207] = 5'b01111; w[102][208] = 5'b01111; w[102][209] = 5'b01111; 
w[103][0] = 5'b01111; w[103][1] = 5'b01111; w[103][2] = 5'b01111; w[103][3] = 5'b01111; w[103][4] = 5'b01111; w[103][5] = 5'b01111; w[103][6] = 5'b01111; w[103][7] = 5'b01111; w[103][8] = 5'b01111; w[103][9] = 5'b01111; w[103][10] = 5'b01111; w[103][11] = 5'b01111; w[103][12] = 5'b01111; w[103][13] = 5'b01111; w[103][14] = 5'b01111; w[103][15] = 5'b01111; w[103][16] = 5'b01111; w[103][17] = 5'b01111; w[103][18] = 5'b01111; w[103][19] = 5'b01111; w[103][20] = 5'b01111; w[103][21] = 5'b01111; w[103][22] = 5'b01111; w[103][23] = 5'b01111; w[103][24] = 5'b01111; w[103][25] = 5'b01111; w[103][26] = 5'b01111; w[103][27] = 5'b01111; w[103][28] = 5'b01111; w[103][29] = 5'b01111; w[103][30] = 5'b01111; w[103][31] = 5'b00000; w[103][32] = 5'b10000; w[103][33] = 5'b10000; w[103][34] = 5'b10000; w[103][35] = 5'b10000; w[103][36] = 5'b10000; w[103][37] = 5'b10000; w[103][38] = 5'b00000; w[103][39] = 5'b01111; w[103][40] = 5'b01111; w[103][41] = 5'b01111; w[103][42] = 5'b01111; w[103][43] = 5'b01111; w[103][44] = 5'b01111; w[103][45] = 5'b10000; w[103][46] = 5'b10000; w[103][47] = 5'b10000; w[103][48] = 5'b10000; w[103][49] = 5'b10000; w[103][50] = 5'b10000; w[103][51] = 5'b10000; w[103][52] = 5'b10000; w[103][53] = 5'b01111; w[103][54] = 5'b01111; w[103][55] = 5'b01111; w[103][56] = 5'b01111; w[103][57] = 5'b01111; w[103][58] = 5'b01111; w[103][59] = 5'b00000; w[103][60] = 5'b00000; w[103][61] = 5'b01111; w[103][62] = 5'b10000; w[103][63] = 5'b00000; w[103][64] = 5'b01111; w[103][65] = 5'b00000; w[103][66] = 5'b00000; w[103][67] = 5'b01111; w[103][68] = 5'b01111; w[103][69] = 5'b01111; w[103][70] = 5'b01111; w[103][71] = 5'b01111; w[103][72] = 5'b01111; w[103][73] = 5'b00000; w[103][74] = 5'b01111; w[103][75] = 5'b01111; w[103][76] = 5'b10000; w[103][77] = 5'b00000; w[103][78] = 5'b01111; w[103][79] = 5'b01111; w[103][80] = 5'b00000; w[103][81] = 5'b01111; w[103][82] = 5'b01111; w[103][83] = 5'b01111; w[103][84] = 5'b01111; w[103][85] = 5'b01111; w[103][86] = 5'b01111; w[103][87] = 5'b00000; w[103][88] = 5'b01111; w[103][89] = 5'b01111; w[103][90] = 5'b10000; w[103][91] = 5'b10000; w[103][92] = 5'b01111; w[103][93] = 5'b01111; w[103][94] = 5'b01111; w[103][95] = 5'b01111; w[103][96] = 5'b01111; w[103][97] = 5'b01111; w[103][98] = 5'b01111; w[103][99] = 5'b01111; w[103][100] = 5'b01111; w[103][101] = 5'b00000; w[103][102] = 5'b01111; w[103][103] = 5'b00000; w[103][104] = 5'b10000; w[103][105] = 5'b10000; w[103][106] = 5'b01111; w[103][107] = 5'b00000; w[103][108] = 5'b00000; w[103][109] = 5'b01111; w[103][110] = 5'b01111; w[103][111] = 5'b01111; w[103][112] = 5'b01111; w[103][113] = 5'b01111; w[103][114] = 5'b01111; w[103][115] = 5'b00000; w[103][116] = 5'b01111; w[103][117] = 5'b01111; w[103][118] = 5'b10000; w[103][119] = 5'b10000; w[103][120] = 5'b00000; w[103][121] = 5'b00000; w[103][122] = 5'b00000; w[103][123] = 5'b01111; w[103][124] = 5'b01111; w[103][125] = 5'b01111; w[103][126] = 5'b01111; w[103][127] = 5'b01111; w[103][128] = 5'b01111; w[103][129] = 5'b00000; w[103][130] = 5'b01111; w[103][131] = 5'b01111; w[103][132] = 5'b00000; w[103][133] = 5'b10000; w[103][134] = 5'b01111; w[103][135] = 5'b01111; w[103][136] = 5'b00000; w[103][137] = 5'b01111; w[103][138] = 5'b01111; w[103][139] = 5'b01111; w[103][140] = 5'b01111; w[103][141] = 5'b01111; w[103][142] = 5'b01111; w[103][143] = 5'b00000; w[103][144] = 5'b00000; w[103][145] = 5'b01111; w[103][146] = 5'b00000; w[103][147] = 5'b10000; w[103][148] = 5'b01111; w[103][149] = 5'b00000; w[103][150] = 5'b00000; w[103][151] = 5'b01111; w[103][152] = 5'b01111; w[103][153] = 5'b01111; w[103][154] = 5'b01111; w[103][155] = 5'b01111; w[103][156] = 5'b01111; w[103][157] = 5'b00000; w[103][158] = 5'b00000; w[103][159] = 5'b00000; w[103][160] = 5'b10000; w[103][161] = 5'b10000; w[103][162] = 5'b10000; w[103][163] = 5'b00000; w[103][164] = 5'b00000; w[103][165] = 5'b01111; w[103][166] = 5'b01111; w[103][167] = 5'b01111; w[103][168] = 5'b01111; w[103][169] = 5'b01111; w[103][170] = 5'b01111; w[103][171] = 5'b01111; w[103][172] = 5'b00000; w[103][173] = 5'b00000; w[103][174] = 5'b10000; w[103][175] = 5'b10000; w[103][176] = 5'b10000; w[103][177] = 5'b00000; w[103][178] = 5'b01111; w[103][179] = 5'b01111; w[103][180] = 5'b01111; w[103][181] = 5'b01111; w[103][182] = 5'b01111; w[103][183] = 5'b01111; w[103][184] = 5'b01111; w[103][185] = 5'b01111; w[103][186] = 5'b01111; w[103][187] = 5'b01111; w[103][188] = 5'b01111; w[103][189] = 5'b01111; w[103][190] = 5'b01111; w[103][191] = 5'b01111; w[103][192] = 5'b01111; w[103][193] = 5'b01111; w[103][194] = 5'b01111; w[103][195] = 5'b01111; w[103][196] = 5'b01111; w[103][197] = 5'b01111; w[103][198] = 5'b01111; w[103][199] = 5'b01111; w[103][200] = 5'b01111; w[103][201] = 5'b01111; w[103][202] = 5'b01111; w[103][203] = 5'b01111; w[103][204] = 5'b01111; w[103][205] = 5'b01111; w[103][206] = 5'b01111; w[103][207] = 5'b01111; w[103][208] = 5'b01111; w[103][209] = 5'b01111; 
w[104][0] = 5'b10000; w[104][1] = 5'b10000; w[104][2] = 5'b10000; w[104][3] = 5'b10000; w[104][4] = 5'b10000; w[104][5] = 5'b10000; w[104][6] = 5'b10000; w[104][7] = 5'b10000; w[104][8] = 5'b10000; w[104][9] = 5'b10000; w[104][10] = 5'b10000; w[104][11] = 5'b10000; w[104][12] = 5'b10000; w[104][13] = 5'b10000; w[104][14] = 5'b10000; w[104][15] = 5'b10000; w[104][16] = 5'b10000; w[104][17] = 5'b10000; w[104][18] = 5'b10000; w[104][19] = 5'b10000; w[104][20] = 5'b10000; w[104][21] = 5'b10000; w[104][22] = 5'b10000; w[104][23] = 5'b10000; w[104][24] = 5'b10000; w[104][25] = 5'b10000; w[104][26] = 5'b10000; w[104][27] = 5'b10000; w[104][28] = 5'b10000; w[104][29] = 5'b10000; w[104][30] = 5'b00000; w[104][31] = 5'b01111; w[104][32] = 5'b00000; w[104][33] = 5'b01111; w[104][34] = 5'b00000; w[104][35] = 5'b00000; w[104][36] = 5'b00000; w[104][37] = 5'b00000; w[104][38] = 5'b01111; w[104][39] = 5'b00000; w[104][40] = 5'b10000; w[104][41] = 5'b10000; w[104][42] = 5'b10000; w[104][43] = 5'b10000; w[104][44] = 5'b00000; w[104][45] = 5'b00000; w[104][46] = 5'b00000; w[104][47] = 5'b01111; w[104][48] = 5'b00000; w[104][49] = 5'b00000; w[104][50] = 5'b00000; w[104][51] = 5'b00000; w[104][52] = 5'b00000; w[104][53] = 5'b00000; w[104][54] = 5'b10000; w[104][55] = 5'b10000; w[104][56] = 5'b10000; w[104][57] = 5'b10000; w[104][58] = 5'b10000; w[104][59] = 5'b10000; w[104][60] = 5'b10000; w[104][61] = 5'b00000; w[104][62] = 5'b01111; w[104][63] = 5'b01111; w[104][64] = 5'b10000; w[104][65] = 5'b10000; w[104][66] = 5'b10000; w[104][67] = 5'b10000; w[104][68] = 5'b10000; w[104][69] = 5'b10000; w[104][70] = 5'b10000; w[104][71] = 5'b10000; w[104][72] = 5'b10000; w[104][73] = 5'b10000; w[104][74] = 5'b00000; w[104][75] = 5'b00000; w[104][76] = 5'b01111; w[104][77] = 5'b01111; w[104][78] = 5'b10000; w[104][79] = 5'b00000; w[104][80] = 5'b10000; w[104][81] = 5'b10000; w[104][82] = 5'b10000; w[104][83] = 5'b10000; w[104][84] = 5'b10000; w[104][85] = 5'b10000; w[104][86] = 5'b10000; w[104][87] = 5'b10000; w[104][88] = 5'b00000; w[104][89] = 5'b00000; w[104][90] = 5'b01111; w[104][91] = 5'b01111; w[104][92] = 5'b10000; w[104][93] = 5'b00000; w[104][94] = 5'b00000; w[104][95] = 5'b10000; w[104][96] = 5'b10000; w[104][97] = 5'b10000; w[104][98] = 5'b10000; w[104][99] = 5'b10000; w[104][100] = 5'b10000; w[104][101] = 5'b10000; w[104][102] = 5'b00000; w[104][103] = 5'b10000; w[104][104] = 5'b00000; w[104][105] = 5'b01111; w[104][106] = 5'b10000; w[104][107] = 5'b10000; w[104][108] = 5'b10000; w[104][109] = 5'b10000; w[104][110] = 5'b10000; w[104][111] = 5'b10000; w[104][112] = 5'b10000; w[104][113] = 5'b10000; w[104][114] = 5'b10000; w[104][115] = 5'b10000; w[104][116] = 5'b00000; w[104][117] = 5'b10000; w[104][118] = 5'b01111; w[104][119] = 5'b01111; w[104][120] = 5'b10000; w[104][121] = 5'b10000; w[104][122] = 5'b10000; w[104][123] = 5'b10000; w[104][124] = 5'b10000; w[104][125] = 5'b10000; w[104][126] = 5'b10000; w[104][127] = 5'b10000; w[104][128] = 5'b10000; w[104][129] = 5'b10000; w[104][130] = 5'b00000; w[104][131] = 5'b10000; w[104][132] = 5'b01111; w[104][133] = 5'b01111; w[104][134] = 5'b00000; w[104][135] = 5'b00000; w[104][136] = 5'b10000; w[104][137] = 5'b10000; w[104][138] = 5'b10000; w[104][139] = 5'b10000; w[104][140] = 5'b10000; w[104][141] = 5'b10000; w[104][142] = 5'b10000; w[104][143] = 5'b10000; w[104][144] = 5'b10000; w[104][145] = 5'b10000; w[104][146] = 5'b01111; w[104][147] = 5'b01111; w[104][148] = 5'b00000; w[104][149] = 5'b10000; w[104][150] = 5'b10000; w[104][151] = 5'b10000; w[104][152] = 5'b10000; w[104][153] = 5'b10000; w[104][154] = 5'b10000; w[104][155] = 5'b10000; w[104][156] = 5'b10000; w[104][157] = 5'b10000; w[104][158] = 5'b10000; w[104][159] = 5'b10000; w[104][160] = 5'b00000; w[104][161] = 5'b00000; w[104][162] = 5'b00000; w[104][163] = 5'b10000; w[104][164] = 5'b10000; w[104][165] = 5'b10000; w[104][166] = 5'b10000; w[104][167] = 5'b10000; w[104][168] = 5'b10000; w[104][169] = 5'b10000; w[104][170] = 5'b10000; w[104][171] = 5'b00000; w[104][172] = 5'b10000; w[104][173] = 5'b10000; w[104][174] = 5'b00000; w[104][175] = 5'b00000; w[104][176] = 5'b00000; w[104][177] = 5'b10000; w[104][178] = 5'b00000; w[104][179] = 5'b10000; w[104][180] = 5'b10000; w[104][181] = 5'b10000; w[104][182] = 5'b10000; w[104][183] = 5'b10000; w[104][184] = 5'b10000; w[104][185] = 5'b10000; w[104][186] = 5'b10000; w[104][187] = 5'b10000; w[104][188] = 5'b10000; w[104][189] = 5'b10000; w[104][190] = 5'b10000; w[104][191] = 5'b10000; w[104][192] = 5'b10000; w[104][193] = 5'b10000; w[104][194] = 5'b10000; w[104][195] = 5'b10000; w[104][196] = 5'b10000; w[104][197] = 5'b10000; w[104][198] = 5'b10000; w[104][199] = 5'b10000; w[104][200] = 5'b10000; w[104][201] = 5'b10000; w[104][202] = 5'b10000; w[104][203] = 5'b10000; w[104][204] = 5'b10000; w[104][205] = 5'b10000; w[104][206] = 5'b10000; w[104][207] = 5'b10000; w[104][208] = 5'b10000; w[104][209] = 5'b10000; 
w[105][0] = 5'b10000; w[105][1] = 5'b10000; w[105][2] = 5'b10000; w[105][3] = 5'b10000; w[105][4] = 5'b10000; w[105][5] = 5'b10000; w[105][6] = 5'b10000; w[105][7] = 5'b10000; w[105][8] = 5'b10000; w[105][9] = 5'b10000; w[105][10] = 5'b10000; w[105][11] = 5'b10000; w[105][12] = 5'b10000; w[105][13] = 5'b10000; w[105][14] = 5'b10000; w[105][15] = 5'b10000; w[105][16] = 5'b10000; w[105][17] = 5'b10000; w[105][18] = 5'b10000; w[105][19] = 5'b10000; w[105][20] = 5'b10000; w[105][21] = 5'b10000; w[105][22] = 5'b10000; w[105][23] = 5'b10000; w[105][24] = 5'b10000; w[105][25] = 5'b10000; w[105][26] = 5'b10000; w[105][27] = 5'b10000; w[105][28] = 5'b10000; w[105][29] = 5'b10000; w[105][30] = 5'b00000; w[105][31] = 5'b01111; w[105][32] = 5'b00000; w[105][33] = 5'b01111; w[105][34] = 5'b00000; w[105][35] = 5'b00000; w[105][36] = 5'b00000; w[105][37] = 5'b00000; w[105][38] = 5'b01111; w[105][39] = 5'b00000; w[105][40] = 5'b10000; w[105][41] = 5'b10000; w[105][42] = 5'b10000; w[105][43] = 5'b10000; w[105][44] = 5'b00000; w[105][45] = 5'b00000; w[105][46] = 5'b00000; w[105][47] = 5'b01111; w[105][48] = 5'b00000; w[105][49] = 5'b00000; w[105][50] = 5'b00000; w[105][51] = 5'b00000; w[105][52] = 5'b00000; w[105][53] = 5'b00000; w[105][54] = 5'b10000; w[105][55] = 5'b10000; w[105][56] = 5'b10000; w[105][57] = 5'b10000; w[105][58] = 5'b10000; w[105][59] = 5'b10000; w[105][60] = 5'b10000; w[105][61] = 5'b00000; w[105][62] = 5'b01111; w[105][63] = 5'b01111; w[105][64] = 5'b10000; w[105][65] = 5'b10000; w[105][66] = 5'b10000; w[105][67] = 5'b10000; w[105][68] = 5'b10000; w[105][69] = 5'b10000; w[105][70] = 5'b10000; w[105][71] = 5'b10000; w[105][72] = 5'b10000; w[105][73] = 5'b10000; w[105][74] = 5'b00000; w[105][75] = 5'b00000; w[105][76] = 5'b01111; w[105][77] = 5'b01111; w[105][78] = 5'b10000; w[105][79] = 5'b00000; w[105][80] = 5'b10000; w[105][81] = 5'b10000; w[105][82] = 5'b10000; w[105][83] = 5'b10000; w[105][84] = 5'b10000; w[105][85] = 5'b10000; w[105][86] = 5'b10000; w[105][87] = 5'b10000; w[105][88] = 5'b00000; w[105][89] = 5'b00000; w[105][90] = 5'b01111; w[105][91] = 5'b01111; w[105][92] = 5'b10000; w[105][93] = 5'b00000; w[105][94] = 5'b00000; w[105][95] = 5'b10000; w[105][96] = 5'b10000; w[105][97] = 5'b10000; w[105][98] = 5'b10000; w[105][99] = 5'b10000; w[105][100] = 5'b10000; w[105][101] = 5'b10000; w[105][102] = 5'b00000; w[105][103] = 5'b10000; w[105][104] = 5'b01111; w[105][105] = 5'b00000; w[105][106] = 5'b10000; w[105][107] = 5'b10000; w[105][108] = 5'b10000; w[105][109] = 5'b10000; w[105][110] = 5'b10000; w[105][111] = 5'b10000; w[105][112] = 5'b10000; w[105][113] = 5'b10000; w[105][114] = 5'b10000; w[105][115] = 5'b10000; w[105][116] = 5'b00000; w[105][117] = 5'b10000; w[105][118] = 5'b01111; w[105][119] = 5'b01111; w[105][120] = 5'b10000; w[105][121] = 5'b10000; w[105][122] = 5'b10000; w[105][123] = 5'b10000; w[105][124] = 5'b10000; w[105][125] = 5'b10000; w[105][126] = 5'b10000; w[105][127] = 5'b10000; w[105][128] = 5'b10000; w[105][129] = 5'b10000; w[105][130] = 5'b00000; w[105][131] = 5'b10000; w[105][132] = 5'b01111; w[105][133] = 5'b01111; w[105][134] = 5'b00000; w[105][135] = 5'b00000; w[105][136] = 5'b10000; w[105][137] = 5'b10000; w[105][138] = 5'b10000; w[105][139] = 5'b10000; w[105][140] = 5'b10000; w[105][141] = 5'b10000; w[105][142] = 5'b10000; w[105][143] = 5'b10000; w[105][144] = 5'b10000; w[105][145] = 5'b10000; w[105][146] = 5'b01111; w[105][147] = 5'b01111; w[105][148] = 5'b00000; w[105][149] = 5'b10000; w[105][150] = 5'b10000; w[105][151] = 5'b10000; w[105][152] = 5'b10000; w[105][153] = 5'b10000; w[105][154] = 5'b10000; w[105][155] = 5'b10000; w[105][156] = 5'b10000; w[105][157] = 5'b10000; w[105][158] = 5'b10000; w[105][159] = 5'b10000; w[105][160] = 5'b00000; w[105][161] = 5'b00000; w[105][162] = 5'b00000; w[105][163] = 5'b10000; w[105][164] = 5'b10000; w[105][165] = 5'b10000; w[105][166] = 5'b10000; w[105][167] = 5'b10000; w[105][168] = 5'b10000; w[105][169] = 5'b10000; w[105][170] = 5'b10000; w[105][171] = 5'b00000; w[105][172] = 5'b10000; w[105][173] = 5'b10000; w[105][174] = 5'b00000; w[105][175] = 5'b00000; w[105][176] = 5'b00000; w[105][177] = 5'b10000; w[105][178] = 5'b00000; w[105][179] = 5'b10000; w[105][180] = 5'b10000; w[105][181] = 5'b10000; w[105][182] = 5'b10000; w[105][183] = 5'b10000; w[105][184] = 5'b10000; w[105][185] = 5'b10000; w[105][186] = 5'b10000; w[105][187] = 5'b10000; w[105][188] = 5'b10000; w[105][189] = 5'b10000; w[105][190] = 5'b10000; w[105][191] = 5'b10000; w[105][192] = 5'b10000; w[105][193] = 5'b10000; w[105][194] = 5'b10000; w[105][195] = 5'b10000; w[105][196] = 5'b10000; w[105][197] = 5'b10000; w[105][198] = 5'b10000; w[105][199] = 5'b10000; w[105][200] = 5'b10000; w[105][201] = 5'b10000; w[105][202] = 5'b10000; w[105][203] = 5'b10000; w[105][204] = 5'b10000; w[105][205] = 5'b10000; w[105][206] = 5'b10000; w[105][207] = 5'b10000; w[105][208] = 5'b10000; w[105][209] = 5'b10000; 
w[106][0] = 5'b01111; w[106][1] = 5'b01111; w[106][2] = 5'b01111; w[106][3] = 5'b01111; w[106][4] = 5'b01111; w[106][5] = 5'b01111; w[106][6] = 5'b01111; w[106][7] = 5'b01111; w[106][8] = 5'b01111; w[106][9] = 5'b01111; w[106][10] = 5'b01111; w[106][11] = 5'b01111; w[106][12] = 5'b01111; w[106][13] = 5'b01111; w[106][14] = 5'b01111; w[106][15] = 5'b01111; w[106][16] = 5'b01111; w[106][17] = 5'b01111; w[106][18] = 5'b01111; w[106][19] = 5'b01111; w[106][20] = 5'b01111; w[106][21] = 5'b01111; w[106][22] = 5'b01111; w[106][23] = 5'b01111; w[106][24] = 5'b01111; w[106][25] = 5'b01111; w[106][26] = 5'b01111; w[106][27] = 5'b01111; w[106][28] = 5'b01111; w[106][29] = 5'b01111; w[106][30] = 5'b00000; w[106][31] = 5'b10000; w[106][32] = 5'b00000; w[106][33] = 5'b10000; w[106][34] = 5'b00000; w[106][35] = 5'b00000; w[106][36] = 5'b00000; w[106][37] = 5'b00000; w[106][38] = 5'b10000; w[106][39] = 5'b00000; w[106][40] = 5'b01111; w[106][41] = 5'b01111; w[106][42] = 5'b01111; w[106][43] = 5'b01111; w[106][44] = 5'b00000; w[106][45] = 5'b00000; w[106][46] = 5'b00000; w[106][47] = 5'b10000; w[106][48] = 5'b00000; w[106][49] = 5'b00000; w[106][50] = 5'b00000; w[106][51] = 5'b00000; w[106][52] = 5'b00000; w[106][53] = 5'b00000; w[106][54] = 5'b01111; w[106][55] = 5'b01111; w[106][56] = 5'b01111; w[106][57] = 5'b01111; w[106][58] = 5'b01111; w[106][59] = 5'b01111; w[106][60] = 5'b01111; w[106][61] = 5'b00000; w[106][62] = 5'b10000; w[106][63] = 5'b10000; w[106][64] = 5'b01111; w[106][65] = 5'b01111; w[106][66] = 5'b01111; w[106][67] = 5'b01111; w[106][68] = 5'b01111; w[106][69] = 5'b01111; w[106][70] = 5'b01111; w[106][71] = 5'b01111; w[106][72] = 5'b01111; w[106][73] = 5'b01111; w[106][74] = 5'b00000; w[106][75] = 5'b00000; w[106][76] = 5'b10000; w[106][77] = 5'b10000; w[106][78] = 5'b01111; w[106][79] = 5'b00000; w[106][80] = 5'b01111; w[106][81] = 5'b01111; w[106][82] = 5'b01111; w[106][83] = 5'b01111; w[106][84] = 5'b01111; w[106][85] = 5'b01111; w[106][86] = 5'b01111; w[106][87] = 5'b01111; w[106][88] = 5'b00000; w[106][89] = 5'b00000; w[106][90] = 5'b10000; w[106][91] = 5'b10000; w[106][92] = 5'b01111; w[106][93] = 5'b00000; w[106][94] = 5'b00000; w[106][95] = 5'b01111; w[106][96] = 5'b01111; w[106][97] = 5'b01111; w[106][98] = 5'b01111; w[106][99] = 5'b01111; w[106][100] = 5'b01111; w[106][101] = 5'b01111; w[106][102] = 5'b00000; w[106][103] = 5'b01111; w[106][104] = 5'b10000; w[106][105] = 5'b10000; w[106][106] = 5'b00000; w[106][107] = 5'b01111; w[106][108] = 5'b01111; w[106][109] = 5'b01111; w[106][110] = 5'b01111; w[106][111] = 5'b01111; w[106][112] = 5'b01111; w[106][113] = 5'b01111; w[106][114] = 5'b01111; w[106][115] = 5'b01111; w[106][116] = 5'b00000; w[106][117] = 5'b01111; w[106][118] = 5'b10000; w[106][119] = 5'b10000; w[106][120] = 5'b01111; w[106][121] = 5'b01111; w[106][122] = 5'b01111; w[106][123] = 5'b01111; w[106][124] = 5'b01111; w[106][125] = 5'b01111; w[106][126] = 5'b01111; w[106][127] = 5'b01111; w[106][128] = 5'b01111; w[106][129] = 5'b01111; w[106][130] = 5'b00000; w[106][131] = 5'b01111; w[106][132] = 5'b10000; w[106][133] = 5'b10000; w[106][134] = 5'b00000; w[106][135] = 5'b00000; w[106][136] = 5'b01111; w[106][137] = 5'b01111; w[106][138] = 5'b01111; w[106][139] = 5'b01111; w[106][140] = 5'b01111; w[106][141] = 5'b01111; w[106][142] = 5'b01111; w[106][143] = 5'b01111; w[106][144] = 5'b01111; w[106][145] = 5'b01111; w[106][146] = 5'b10000; w[106][147] = 5'b10000; w[106][148] = 5'b00000; w[106][149] = 5'b01111; w[106][150] = 5'b01111; w[106][151] = 5'b01111; w[106][152] = 5'b01111; w[106][153] = 5'b01111; w[106][154] = 5'b01111; w[106][155] = 5'b01111; w[106][156] = 5'b01111; w[106][157] = 5'b01111; w[106][158] = 5'b01111; w[106][159] = 5'b01111; w[106][160] = 5'b00000; w[106][161] = 5'b00000; w[106][162] = 5'b00000; w[106][163] = 5'b01111; w[106][164] = 5'b01111; w[106][165] = 5'b01111; w[106][166] = 5'b01111; w[106][167] = 5'b01111; w[106][168] = 5'b01111; w[106][169] = 5'b01111; w[106][170] = 5'b01111; w[106][171] = 5'b00000; w[106][172] = 5'b01111; w[106][173] = 5'b01111; w[106][174] = 5'b00000; w[106][175] = 5'b00000; w[106][176] = 5'b00000; w[106][177] = 5'b01111; w[106][178] = 5'b00000; w[106][179] = 5'b01111; w[106][180] = 5'b01111; w[106][181] = 5'b01111; w[106][182] = 5'b01111; w[106][183] = 5'b01111; w[106][184] = 5'b01111; w[106][185] = 5'b01111; w[106][186] = 5'b01111; w[106][187] = 5'b01111; w[106][188] = 5'b01111; w[106][189] = 5'b01111; w[106][190] = 5'b01111; w[106][191] = 5'b01111; w[106][192] = 5'b01111; w[106][193] = 5'b01111; w[106][194] = 5'b01111; w[106][195] = 5'b01111; w[106][196] = 5'b01111; w[106][197] = 5'b01111; w[106][198] = 5'b01111; w[106][199] = 5'b01111; w[106][200] = 5'b01111; w[106][201] = 5'b01111; w[106][202] = 5'b01111; w[106][203] = 5'b01111; w[106][204] = 5'b01111; w[106][205] = 5'b01111; w[106][206] = 5'b01111; w[106][207] = 5'b01111; w[106][208] = 5'b01111; w[106][209] = 5'b01111; 
w[107][0] = 5'b00000; w[107][1] = 5'b00000; w[107][2] = 5'b00000; w[107][3] = 5'b00000; w[107][4] = 5'b00000; w[107][5] = 5'b00000; w[107][6] = 5'b00000; w[107][7] = 5'b00000; w[107][8] = 5'b00000; w[107][9] = 5'b00000; w[107][10] = 5'b00000; w[107][11] = 5'b00000; w[107][12] = 5'b00000; w[107][13] = 5'b00000; w[107][14] = 5'b00000; w[107][15] = 5'b00000; w[107][16] = 5'b00000; w[107][17] = 5'b00000; w[107][18] = 5'b00000; w[107][19] = 5'b00000; w[107][20] = 5'b00000; w[107][21] = 5'b00000; w[107][22] = 5'b00000; w[107][23] = 5'b00000; w[107][24] = 5'b00000; w[107][25] = 5'b00000; w[107][26] = 5'b00000; w[107][27] = 5'b00000; w[107][28] = 5'b00000; w[107][29] = 5'b00000; w[107][30] = 5'b10000; w[107][31] = 5'b00000; w[107][32] = 5'b01111; w[107][33] = 5'b00000; w[107][34] = 5'b10000; w[107][35] = 5'b10000; w[107][36] = 5'b10000; w[107][37] = 5'b01111; w[107][38] = 5'b00000; w[107][39] = 5'b10000; w[107][40] = 5'b00000; w[107][41] = 5'b00000; w[107][42] = 5'b00000; w[107][43] = 5'b00000; w[107][44] = 5'b10000; w[107][45] = 5'b01111; w[107][46] = 5'b01111; w[107][47] = 5'b00000; w[107][48] = 5'b10000; w[107][49] = 5'b10000; w[107][50] = 5'b10000; w[107][51] = 5'b01111; w[107][52] = 5'b01111; w[107][53] = 5'b10000; w[107][54] = 5'b00000; w[107][55] = 5'b00000; w[107][56] = 5'b00000; w[107][57] = 5'b00000; w[107][58] = 5'b01111; w[107][59] = 5'b01111; w[107][60] = 5'b01111; w[107][61] = 5'b01111; w[107][62] = 5'b10000; w[107][63] = 5'b10000; w[107][64] = 5'b00000; w[107][65] = 5'b01111; w[107][66] = 5'b01111; w[107][67] = 5'b01111; w[107][68] = 5'b00000; w[107][69] = 5'b00000; w[107][70] = 5'b00000; w[107][71] = 5'b00000; w[107][72] = 5'b01111; w[107][73] = 5'b01111; w[107][74] = 5'b01111; w[107][75] = 5'b01111; w[107][76] = 5'b10000; w[107][77] = 5'b10000; w[107][78] = 5'b00000; w[107][79] = 5'b01111; w[107][80] = 5'b01111; w[107][81] = 5'b01111; w[107][82] = 5'b00000; w[107][83] = 5'b00000; w[107][84] = 5'b00000; w[107][85] = 5'b00000; w[107][86] = 5'b01111; w[107][87] = 5'b01111; w[107][88] = 5'b01111; w[107][89] = 5'b01111; w[107][90] = 5'b10000; w[107][91] = 5'b10000; w[107][92] = 5'b00000; w[107][93] = 5'b01111; w[107][94] = 5'b01111; w[107][95] = 5'b00000; w[107][96] = 5'b00000; w[107][97] = 5'b00000; w[107][98] = 5'b00000; w[107][99] = 5'b00000; w[107][100] = 5'b01111; w[107][101] = 5'b01111; w[107][102] = 5'b01111; w[107][103] = 5'b00000; w[107][104] = 5'b10000; w[107][105] = 5'b10000; w[107][106] = 5'b01111; w[107][107] = 5'b00000; w[107][108] = 5'b01111; w[107][109] = 5'b01111; w[107][110] = 5'b00000; w[107][111] = 5'b00000; w[107][112] = 5'b00000; w[107][113] = 5'b00000; w[107][114] = 5'b01111; w[107][115] = 5'b01111; w[107][116] = 5'b01111; w[107][117] = 5'b00000; w[107][118] = 5'b10000; w[107][119] = 5'b10000; w[107][120] = 5'b01111; w[107][121] = 5'b01111; w[107][122] = 5'b01111; w[107][123] = 5'b01111; w[107][124] = 5'b00000; w[107][125] = 5'b00000; w[107][126] = 5'b00000; w[107][127] = 5'b00000; w[107][128] = 5'b01111; w[107][129] = 5'b01111; w[107][130] = 5'b01111; w[107][131] = 5'b00000; w[107][132] = 5'b10000; w[107][133] = 5'b10000; w[107][134] = 5'b01111; w[107][135] = 5'b01111; w[107][136] = 5'b01111; w[107][137] = 5'b01111; w[107][138] = 5'b00000; w[107][139] = 5'b00000; w[107][140] = 5'b00000; w[107][141] = 5'b00000; w[107][142] = 5'b01111; w[107][143] = 5'b01111; w[107][144] = 5'b01111; w[107][145] = 5'b00000; w[107][146] = 5'b10000; w[107][147] = 5'b10000; w[107][148] = 5'b01111; w[107][149] = 5'b01111; w[107][150] = 5'b01111; w[107][151] = 5'b01111; w[107][152] = 5'b00000; w[107][153] = 5'b00000; w[107][154] = 5'b00000; w[107][155] = 5'b00000; w[107][156] = 5'b00000; w[107][157] = 5'b01111; w[107][158] = 5'b01111; w[107][159] = 5'b00000; w[107][160] = 5'b10000; w[107][161] = 5'b10000; w[107][162] = 5'b01111; w[107][163] = 5'b01111; w[107][164] = 5'b01111; w[107][165] = 5'b00000; w[107][166] = 5'b00000; w[107][167] = 5'b00000; w[107][168] = 5'b00000; w[107][169] = 5'b00000; w[107][170] = 5'b00000; w[107][171] = 5'b01111; w[107][172] = 5'b01111; w[107][173] = 5'b00000; w[107][174] = 5'b10000; w[107][175] = 5'b10000; w[107][176] = 5'b01111; w[107][177] = 5'b01111; w[107][178] = 5'b01111; w[107][179] = 5'b00000; w[107][180] = 5'b00000; w[107][181] = 5'b00000; w[107][182] = 5'b00000; w[107][183] = 5'b00000; w[107][184] = 5'b00000; w[107][185] = 5'b00000; w[107][186] = 5'b00000; w[107][187] = 5'b00000; w[107][188] = 5'b00000; w[107][189] = 5'b00000; w[107][190] = 5'b00000; w[107][191] = 5'b00000; w[107][192] = 5'b00000; w[107][193] = 5'b00000; w[107][194] = 5'b00000; w[107][195] = 5'b00000; w[107][196] = 5'b00000; w[107][197] = 5'b00000; w[107][198] = 5'b00000; w[107][199] = 5'b00000; w[107][200] = 5'b00000; w[107][201] = 5'b00000; w[107][202] = 5'b00000; w[107][203] = 5'b00000; w[107][204] = 5'b00000; w[107][205] = 5'b00000; w[107][206] = 5'b00000; w[107][207] = 5'b00000; w[107][208] = 5'b00000; w[107][209] = 5'b00000; 
w[108][0] = 5'b00000; w[108][1] = 5'b00000; w[108][2] = 5'b00000; w[108][3] = 5'b00000; w[108][4] = 5'b00000; w[108][5] = 5'b00000; w[108][6] = 5'b00000; w[108][7] = 5'b00000; w[108][8] = 5'b00000; w[108][9] = 5'b00000; w[108][10] = 5'b00000; w[108][11] = 5'b00000; w[108][12] = 5'b00000; w[108][13] = 5'b00000; w[108][14] = 5'b00000; w[108][15] = 5'b00000; w[108][16] = 5'b00000; w[108][17] = 5'b00000; w[108][18] = 5'b00000; w[108][19] = 5'b00000; w[108][20] = 5'b00000; w[108][21] = 5'b00000; w[108][22] = 5'b00000; w[108][23] = 5'b00000; w[108][24] = 5'b00000; w[108][25] = 5'b00000; w[108][26] = 5'b00000; w[108][27] = 5'b00000; w[108][28] = 5'b00000; w[108][29] = 5'b00000; w[108][30] = 5'b10000; w[108][31] = 5'b00000; w[108][32] = 5'b01111; w[108][33] = 5'b00000; w[108][34] = 5'b10000; w[108][35] = 5'b10000; w[108][36] = 5'b10000; w[108][37] = 5'b01111; w[108][38] = 5'b00000; w[108][39] = 5'b10000; w[108][40] = 5'b00000; w[108][41] = 5'b00000; w[108][42] = 5'b00000; w[108][43] = 5'b00000; w[108][44] = 5'b10000; w[108][45] = 5'b01111; w[108][46] = 5'b01111; w[108][47] = 5'b00000; w[108][48] = 5'b10000; w[108][49] = 5'b10000; w[108][50] = 5'b10000; w[108][51] = 5'b01111; w[108][52] = 5'b01111; w[108][53] = 5'b10000; w[108][54] = 5'b00000; w[108][55] = 5'b00000; w[108][56] = 5'b00000; w[108][57] = 5'b00000; w[108][58] = 5'b01111; w[108][59] = 5'b01111; w[108][60] = 5'b01111; w[108][61] = 5'b01111; w[108][62] = 5'b10000; w[108][63] = 5'b10000; w[108][64] = 5'b00000; w[108][65] = 5'b01111; w[108][66] = 5'b01111; w[108][67] = 5'b01111; w[108][68] = 5'b00000; w[108][69] = 5'b00000; w[108][70] = 5'b00000; w[108][71] = 5'b00000; w[108][72] = 5'b01111; w[108][73] = 5'b01111; w[108][74] = 5'b01111; w[108][75] = 5'b01111; w[108][76] = 5'b10000; w[108][77] = 5'b10000; w[108][78] = 5'b00000; w[108][79] = 5'b01111; w[108][80] = 5'b01111; w[108][81] = 5'b01111; w[108][82] = 5'b00000; w[108][83] = 5'b00000; w[108][84] = 5'b00000; w[108][85] = 5'b00000; w[108][86] = 5'b01111; w[108][87] = 5'b01111; w[108][88] = 5'b01111; w[108][89] = 5'b01111; w[108][90] = 5'b10000; w[108][91] = 5'b10000; w[108][92] = 5'b00000; w[108][93] = 5'b01111; w[108][94] = 5'b01111; w[108][95] = 5'b00000; w[108][96] = 5'b00000; w[108][97] = 5'b00000; w[108][98] = 5'b00000; w[108][99] = 5'b00000; w[108][100] = 5'b01111; w[108][101] = 5'b01111; w[108][102] = 5'b01111; w[108][103] = 5'b00000; w[108][104] = 5'b10000; w[108][105] = 5'b10000; w[108][106] = 5'b01111; w[108][107] = 5'b01111; w[108][108] = 5'b00000; w[108][109] = 5'b01111; w[108][110] = 5'b00000; w[108][111] = 5'b00000; w[108][112] = 5'b00000; w[108][113] = 5'b00000; w[108][114] = 5'b01111; w[108][115] = 5'b01111; w[108][116] = 5'b01111; w[108][117] = 5'b00000; w[108][118] = 5'b10000; w[108][119] = 5'b10000; w[108][120] = 5'b01111; w[108][121] = 5'b01111; w[108][122] = 5'b01111; w[108][123] = 5'b01111; w[108][124] = 5'b00000; w[108][125] = 5'b00000; w[108][126] = 5'b00000; w[108][127] = 5'b00000; w[108][128] = 5'b01111; w[108][129] = 5'b01111; w[108][130] = 5'b01111; w[108][131] = 5'b00000; w[108][132] = 5'b10000; w[108][133] = 5'b10000; w[108][134] = 5'b01111; w[108][135] = 5'b01111; w[108][136] = 5'b01111; w[108][137] = 5'b01111; w[108][138] = 5'b00000; w[108][139] = 5'b00000; w[108][140] = 5'b00000; w[108][141] = 5'b00000; w[108][142] = 5'b01111; w[108][143] = 5'b01111; w[108][144] = 5'b01111; w[108][145] = 5'b00000; w[108][146] = 5'b10000; w[108][147] = 5'b10000; w[108][148] = 5'b01111; w[108][149] = 5'b01111; w[108][150] = 5'b01111; w[108][151] = 5'b01111; w[108][152] = 5'b00000; w[108][153] = 5'b00000; w[108][154] = 5'b00000; w[108][155] = 5'b00000; w[108][156] = 5'b00000; w[108][157] = 5'b01111; w[108][158] = 5'b01111; w[108][159] = 5'b00000; w[108][160] = 5'b10000; w[108][161] = 5'b10000; w[108][162] = 5'b01111; w[108][163] = 5'b01111; w[108][164] = 5'b01111; w[108][165] = 5'b00000; w[108][166] = 5'b00000; w[108][167] = 5'b00000; w[108][168] = 5'b00000; w[108][169] = 5'b00000; w[108][170] = 5'b00000; w[108][171] = 5'b01111; w[108][172] = 5'b01111; w[108][173] = 5'b00000; w[108][174] = 5'b10000; w[108][175] = 5'b10000; w[108][176] = 5'b01111; w[108][177] = 5'b01111; w[108][178] = 5'b01111; w[108][179] = 5'b00000; w[108][180] = 5'b00000; w[108][181] = 5'b00000; w[108][182] = 5'b00000; w[108][183] = 5'b00000; w[108][184] = 5'b00000; w[108][185] = 5'b00000; w[108][186] = 5'b00000; w[108][187] = 5'b00000; w[108][188] = 5'b00000; w[108][189] = 5'b00000; w[108][190] = 5'b00000; w[108][191] = 5'b00000; w[108][192] = 5'b00000; w[108][193] = 5'b00000; w[108][194] = 5'b00000; w[108][195] = 5'b00000; w[108][196] = 5'b00000; w[108][197] = 5'b00000; w[108][198] = 5'b00000; w[108][199] = 5'b00000; w[108][200] = 5'b00000; w[108][201] = 5'b00000; w[108][202] = 5'b00000; w[108][203] = 5'b00000; w[108][204] = 5'b00000; w[108][205] = 5'b00000; w[108][206] = 5'b00000; w[108][207] = 5'b00000; w[108][208] = 5'b00000; w[108][209] = 5'b00000; 
w[109][0] = 5'b01111; w[109][1] = 5'b01111; w[109][2] = 5'b01111; w[109][3] = 5'b01111; w[109][4] = 5'b01111; w[109][5] = 5'b01111; w[109][6] = 5'b01111; w[109][7] = 5'b01111; w[109][8] = 5'b01111; w[109][9] = 5'b01111; w[109][10] = 5'b01111; w[109][11] = 5'b01111; w[109][12] = 5'b01111; w[109][13] = 5'b01111; w[109][14] = 5'b01111; w[109][15] = 5'b01111; w[109][16] = 5'b01111; w[109][17] = 5'b01111; w[109][18] = 5'b01111; w[109][19] = 5'b01111; w[109][20] = 5'b01111; w[109][21] = 5'b01111; w[109][22] = 5'b01111; w[109][23] = 5'b01111; w[109][24] = 5'b01111; w[109][25] = 5'b01111; w[109][26] = 5'b01111; w[109][27] = 5'b01111; w[109][28] = 5'b01111; w[109][29] = 5'b01111; w[109][30] = 5'b00000; w[109][31] = 5'b10000; w[109][32] = 5'b00000; w[109][33] = 5'b10000; w[109][34] = 5'b00000; w[109][35] = 5'b00000; w[109][36] = 5'b00000; w[109][37] = 5'b00000; w[109][38] = 5'b10000; w[109][39] = 5'b00000; w[109][40] = 5'b01111; w[109][41] = 5'b01111; w[109][42] = 5'b01111; w[109][43] = 5'b01111; w[109][44] = 5'b00000; w[109][45] = 5'b00000; w[109][46] = 5'b00000; w[109][47] = 5'b10000; w[109][48] = 5'b00000; w[109][49] = 5'b00000; w[109][50] = 5'b00000; w[109][51] = 5'b00000; w[109][52] = 5'b00000; w[109][53] = 5'b00000; w[109][54] = 5'b01111; w[109][55] = 5'b01111; w[109][56] = 5'b01111; w[109][57] = 5'b01111; w[109][58] = 5'b01111; w[109][59] = 5'b01111; w[109][60] = 5'b01111; w[109][61] = 5'b00000; w[109][62] = 5'b10000; w[109][63] = 5'b10000; w[109][64] = 5'b01111; w[109][65] = 5'b01111; w[109][66] = 5'b01111; w[109][67] = 5'b01111; w[109][68] = 5'b01111; w[109][69] = 5'b01111; w[109][70] = 5'b01111; w[109][71] = 5'b01111; w[109][72] = 5'b01111; w[109][73] = 5'b01111; w[109][74] = 5'b00000; w[109][75] = 5'b00000; w[109][76] = 5'b10000; w[109][77] = 5'b10000; w[109][78] = 5'b01111; w[109][79] = 5'b00000; w[109][80] = 5'b01111; w[109][81] = 5'b01111; w[109][82] = 5'b01111; w[109][83] = 5'b01111; w[109][84] = 5'b01111; w[109][85] = 5'b01111; w[109][86] = 5'b01111; w[109][87] = 5'b01111; w[109][88] = 5'b00000; w[109][89] = 5'b00000; w[109][90] = 5'b10000; w[109][91] = 5'b10000; w[109][92] = 5'b01111; w[109][93] = 5'b00000; w[109][94] = 5'b00000; w[109][95] = 5'b01111; w[109][96] = 5'b01111; w[109][97] = 5'b01111; w[109][98] = 5'b01111; w[109][99] = 5'b01111; w[109][100] = 5'b01111; w[109][101] = 5'b01111; w[109][102] = 5'b00000; w[109][103] = 5'b01111; w[109][104] = 5'b10000; w[109][105] = 5'b10000; w[109][106] = 5'b01111; w[109][107] = 5'b01111; w[109][108] = 5'b01111; w[109][109] = 5'b00000; w[109][110] = 5'b01111; w[109][111] = 5'b01111; w[109][112] = 5'b01111; w[109][113] = 5'b01111; w[109][114] = 5'b01111; w[109][115] = 5'b01111; w[109][116] = 5'b00000; w[109][117] = 5'b01111; w[109][118] = 5'b10000; w[109][119] = 5'b10000; w[109][120] = 5'b01111; w[109][121] = 5'b01111; w[109][122] = 5'b01111; w[109][123] = 5'b01111; w[109][124] = 5'b01111; w[109][125] = 5'b01111; w[109][126] = 5'b01111; w[109][127] = 5'b01111; w[109][128] = 5'b01111; w[109][129] = 5'b01111; w[109][130] = 5'b00000; w[109][131] = 5'b01111; w[109][132] = 5'b10000; w[109][133] = 5'b10000; w[109][134] = 5'b00000; w[109][135] = 5'b00000; w[109][136] = 5'b01111; w[109][137] = 5'b01111; w[109][138] = 5'b01111; w[109][139] = 5'b01111; w[109][140] = 5'b01111; w[109][141] = 5'b01111; w[109][142] = 5'b01111; w[109][143] = 5'b01111; w[109][144] = 5'b01111; w[109][145] = 5'b01111; w[109][146] = 5'b10000; w[109][147] = 5'b10000; w[109][148] = 5'b00000; w[109][149] = 5'b01111; w[109][150] = 5'b01111; w[109][151] = 5'b01111; w[109][152] = 5'b01111; w[109][153] = 5'b01111; w[109][154] = 5'b01111; w[109][155] = 5'b01111; w[109][156] = 5'b01111; w[109][157] = 5'b01111; w[109][158] = 5'b01111; w[109][159] = 5'b01111; w[109][160] = 5'b00000; w[109][161] = 5'b00000; w[109][162] = 5'b00000; w[109][163] = 5'b01111; w[109][164] = 5'b01111; w[109][165] = 5'b01111; w[109][166] = 5'b01111; w[109][167] = 5'b01111; w[109][168] = 5'b01111; w[109][169] = 5'b01111; w[109][170] = 5'b01111; w[109][171] = 5'b00000; w[109][172] = 5'b01111; w[109][173] = 5'b01111; w[109][174] = 5'b00000; w[109][175] = 5'b00000; w[109][176] = 5'b00000; w[109][177] = 5'b01111; w[109][178] = 5'b00000; w[109][179] = 5'b01111; w[109][180] = 5'b01111; w[109][181] = 5'b01111; w[109][182] = 5'b01111; w[109][183] = 5'b01111; w[109][184] = 5'b01111; w[109][185] = 5'b01111; w[109][186] = 5'b01111; w[109][187] = 5'b01111; w[109][188] = 5'b01111; w[109][189] = 5'b01111; w[109][190] = 5'b01111; w[109][191] = 5'b01111; w[109][192] = 5'b01111; w[109][193] = 5'b01111; w[109][194] = 5'b01111; w[109][195] = 5'b01111; w[109][196] = 5'b01111; w[109][197] = 5'b01111; w[109][198] = 5'b01111; w[109][199] = 5'b01111; w[109][200] = 5'b01111; w[109][201] = 5'b01111; w[109][202] = 5'b01111; w[109][203] = 5'b01111; w[109][204] = 5'b01111; w[109][205] = 5'b01111; w[109][206] = 5'b01111; w[109][207] = 5'b01111; w[109][208] = 5'b01111; w[109][209] = 5'b01111; 
w[110][0] = 5'b01111; w[110][1] = 5'b01111; w[110][2] = 5'b01111; w[110][3] = 5'b01111; w[110][4] = 5'b01111; w[110][5] = 5'b01111; w[110][6] = 5'b01111; w[110][7] = 5'b01111; w[110][8] = 5'b01111; w[110][9] = 5'b01111; w[110][10] = 5'b01111; w[110][11] = 5'b01111; w[110][12] = 5'b01111; w[110][13] = 5'b01111; w[110][14] = 5'b01111; w[110][15] = 5'b01111; w[110][16] = 5'b01111; w[110][17] = 5'b01111; w[110][18] = 5'b01111; w[110][19] = 5'b01111; w[110][20] = 5'b01111; w[110][21] = 5'b01111; w[110][22] = 5'b01111; w[110][23] = 5'b01111; w[110][24] = 5'b01111; w[110][25] = 5'b01111; w[110][26] = 5'b01111; w[110][27] = 5'b01111; w[110][28] = 5'b01111; w[110][29] = 5'b01111; w[110][30] = 5'b01111; w[110][31] = 5'b00000; w[110][32] = 5'b10000; w[110][33] = 5'b10000; w[110][34] = 5'b10000; w[110][35] = 5'b10000; w[110][36] = 5'b10000; w[110][37] = 5'b10000; w[110][38] = 5'b00000; w[110][39] = 5'b01111; w[110][40] = 5'b01111; w[110][41] = 5'b01111; w[110][42] = 5'b01111; w[110][43] = 5'b01111; w[110][44] = 5'b01111; w[110][45] = 5'b10000; w[110][46] = 5'b10000; w[110][47] = 5'b10000; w[110][48] = 5'b10000; w[110][49] = 5'b10000; w[110][50] = 5'b10000; w[110][51] = 5'b10000; w[110][52] = 5'b10000; w[110][53] = 5'b01111; w[110][54] = 5'b01111; w[110][55] = 5'b01111; w[110][56] = 5'b01111; w[110][57] = 5'b01111; w[110][58] = 5'b01111; w[110][59] = 5'b00000; w[110][60] = 5'b00000; w[110][61] = 5'b01111; w[110][62] = 5'b10000; w[110][63] = 5'b00000; w[110][64] = 5'b01111; w[110][65] = 5'b00000; w[110][66] = 5'b00000; w[110][67] = 5'b01111; w[110][68] = 5'b01111; w[110][69] = 5'b01111; w[110][70] = 5'b01111; w[110][71] = 5'b01111; w[110][72] = 5'b01111; w[110][73] = 5'b00000; w[110][74] = 5'b01111; w[110][75] = 5'b01111; w[110][76] = 5'b10000; w[110][77] = 5'b00000; w[110][78] = 5'b01111; w[110][79] = 5'b01111; w[110][80] = 5'b00000; w[110][81] = 5'b01111; w[110][82] = 5'b01111; w[110][83] = 5'b01111; w[110][84] = 5'b01111; w[110][85] = 5'b01111; w[110][86] = 5'b01111; w[110][87] = 5'b00000; w[110][88] = 5'b01111; w[110][89] = 5'b01111; w[110][90] = 5'b10000; w[110][91] = 5'b10000; w[110][92] = 5'b01111; w[110][93] = 5'b01111; w[110][94] = 5'b01111; w[110][95] = 5'b01111; w[110][96] = 5'b01111; w[110][97] = 5'b01111; w[110][98] = 5'b01111; w[110][99] = 5'b01111; w[110][100] = 5'b01111; w[110][101] = 5'b00000; w[110][102] = 5'b01111; w[110][103] = 5'b01111; w[110][104] = 5'b10000; w[110][105] = 5'b10000; w[110][106] = 5'b01111; w[110][107] = 5'b00000; w[110][108] = 5'b00000; w[110][109] = 5'b01111; w[110][110] = 5'b00000; w[110][111] = 5'b01111; w[110][112] = 5'b01111; w[110][113] = 5'b01111; w[110][114] = 5'b01111; w[110][115] = 5'b00000; w[110][116] = 5'b01111; w[110][117] = 5'b01111; w[110][118] = 5'b10000; w[110][119] = 5'b10000; w[110][120] = 5'b00000; w[110][121] = 5'b00000; w[110][122] = 5'b00000; w[110][123] = 5'b01111; w[110][124] = 5'b01111; w[110][125] = 5'b01111; w[110][126] = 5'b01111; w[110][127] = 5'b01111; w[110][128] = 5'b01111; w[110][129] = 5'b00000; w[110][130] = 5'b01111; w[110][131] = 5'b01111; w[110][132] = 5'b00000; w[110][133] = 5'b10000; w[110][134] = 5'b01111; w[110][135] = 5'b01111; w[110][136] = 5'b00000; w[110][137] = 5'b01111; w[110][138] = 5'b01111; w[110][139] = 5'b01111; w[110][140] = 5'b01111; w[110][141] = 5'b01111; w[110][142] = 5'b01111; w[110][143] = 5'b00000; w[110][144] = 5'b00000; w[110][145] = 5'b01111; w[110][146] = 5'b00000; w[110][147] = 5'b10000; w[110][148] = 5'b01111; w[110][149] = 5'b00000; w[110][150] = 5'b00000; w[110][151] = 5'b01111; w[110][152] = 5'b01111; w[110][153] = 5'b01111; w[110][154] = 5'b01111; w[110][155] = 5'b01111; w[110][156] = 5'b01111; w[110][157] = 5'b00000; w[110][158] = 5'b00000; w[110][159] = 5'b00000; w[110][160] = 5'b10000; w[110][161] = 5'b10000; w[110][162] = 5'b10000; w[110][163] = 5'b00000; w[110][164] = 5'b00000; w[110][165] = 5'b01111; w[110][166] = 5'b01111; w[110][167] = 5'b01111; w[110][168] = 5'b01111; w[110][169] = 5'b01111; w[110][170] = 5'b01111; w[110][171] = 5'b01111; w[110][172] = 5'b00000; w[110][173] = 5'b00000; w[110][174] = 5'b10000; w[110][175] = 5'b10000; w[110][176] = 5'b10000; w[110][177] = 5'b00000; w[110][178] = 5'b01111; w[110][179] = 5'b01111; w[110][180] = 5'b01111; w[110][181] = 5'b01111; w[110][182] = 5'b01111; w[110][183] = 5'b01111; w[110][184] = 5'b01111; w[110][185] = 5'b01111; w[110][186] = 5'b01111; w[110][187] = 5'b01111; w[110][188] = 5'b01111; w[110][189] = 5'b01111; w[110][190] = 5'b01111; w[110][191] = 5'b01111; w[110][192] = 5'b01111; w[110][193] = 5'b01111; w[110][194] = 5'b01111; w[110][195] = 5'b01111; w[110][196] = 5'b01111; w[110][197] = 5'b01111; w[110][198] = 5'b01111; w[110][199] = 5'b01111; w[110][200] = 5'b01111; w[110][201] = 5'b01111; w[110][202] = 5'b01111; w[110][203] = 5'b01111; w[110][204] = 5'b01111; w[110][205] = 5'b01111; w[110][206] = 5'b01111; w[110][207] = 5'b01111; w[110][208] = 5'b01111; w[110][209] = 5'b01111; 
w[111][0] = 5'b01111; w[111][1] = 5'b01111; w[111][2] = 5'b01111; w[111][3] = 5'b01111; w[111][4] = 5'b01111; w[111][5] = 5'b01111; w[111][6] = 5'b01111; w[111][7] = 5'b01111; w[111][8] = 5'b01111; w[111][9] = 5'b01111; w[111][10] = 5'b01111; w[111][11] = 5'b01111; w[111][12] = 5'b01111; w[111][13] = 5'b01111; w[111][14] = 5'b01111; w[111][15] = 5'b01111; w[111][16] = 5'b01111; w[111][17] = 5'b01111; w[111][18] = 5'b01111; w[111][19] = 5'b01111; w[111][20] = 5'b01111; w[111][21] = 5'b01111; w[111][22] = 5'b01111; w[111][23] = 5'b01111; w[111][24] = 5'b01111; w[111][25] = 5'b01111; w[111][26] = 5'b01111; w[111][27] = 5'b01111; w[111][28] = 5'b01111; w[111][29] = 5'b01111; w[111][30] = 5'b01111; w[111][31] = 5'b00000; w[111][32] = 5'b10000; w[111][33] = 5'b10000; w[111][34] = 5'b10000; w[111][35] = 5'b10000; w[111][36] = 5'b10000; w[111][37] = 5'b10000; w[111][38] = 5'b00000; w[111][39] = 5'b01111; w[111][40] = 5'b01111; w[111][41] = 5'b01111; w[111][42] = 5'b01111; w[111][43] = 5'b01111; w[111][44] = 5'b01111; w[111][45] = 5'b10000; w[111][46] = 5'b10000; w[111][47] = 5'b10000; w[111][48] = 5'b10000; w[111][49] = 5'b10000; w[111][50] = 5'b10000; w[111][51] = 5'b10000; w[111][52] = 5'b10000; w[111][53] = 5'b01111; w[111][54] = 5'b01111; w[111][55] = 5'b01111; w[111][56] = 5'b01111; w[111][57] = 5'b01111; w[111][58] = 5'b01111; w[111][59] = 5'b00000; w[111][60] = 5'b00000; w[111][61] = 5'b01111; w[111][62] = 5'b10000; w[111][63] = 5'b00000; w[111][64] = 5'b01111; w[111][65] = 5'b00000; w[111][66] = 5'b00000; w[111][67] = 5'b01111; w[111][68] = 5'b01111; w[111][69] = 5'b01111; w[111][70] = 5'b01111; w[111][71] = 5'b01111; w[111][72] = 5'b01111; w[111][73] = 5'b00000; w[111][74] = 5'b01111; w[111][75] = 5'b01111; w[111][76] = 5'b10000; w[111][77] = 5'b00000; w[111][78] = 5'b01111; w[111][79] = 5'b01111; w[111][80] = 5'b00000; w[111][81] = 5'b01111; w[111][82] = 5'b01111; w[111][83] = 5'b01111; w[111][84] = 5'b01111; w[111][85] = 5'b01111; w[111][86] = 5'b01111; w[111][87] = 5'b00000; w[111][88] = 5'b01111; w[111][89] = 5'b01111; w[111][90] = 5'b10000; w[111][91] = 5'b10000; w[111][92] = 5'b01111; w[111][93] = 5'b01111; w[111][94] = 5'b01111; w[111][95] = 5'b01111; w[111][96] = 5'b01111; w[111][97] = 5'b01111; w[111][98] = 5'b01111; w[111][99] = 5'b01111; w[111][100] = 5'b01111; w[111][101] = 5'b00000; w[111][102] = 5'b01111; w[111][103] = 5'b01111; w[111][104] = 5'b10000; w[111][105] = 5'b10000; w[111][106] = 5'b01111; w[111][107] = 5'b00000; w[111][108] = 5'b00000; w[111][109] = 5'b01111; w[111][110] = 5'b01111; w[111][111] = 5'b00000; w[111][112] = 5'b01111; w[111][113] = 5'b01111; w[111][114] = 5'b01111; w[111][115] = 5'b00000; w[111][116] = 5'b01111; w[111][117] = 5'b01111; w[111][118] = 5'b10000; w[111][119] = 5'b10000; w[111][120] = 5'b00000; w[111][121] = 5'b00000; w[111][122] = 5'b00000; w[111][123] = 5'b01111; w[111][124] = 5'b01111; w[111][125] = 5'b01111; w[111][126] = 5'b01111; w[111][127] = 5'b01111; w[111][128] = 5'b01111; w[111][129] = 5'b00000; w[111][130] = 5'b01111; w[111][131] = 5'b01111; w[111][132] = 5'b00000; w[111][133] = 5'b10000; w[111][134] = 5'b01111; w[111][135] = 5'b01111; w[111][136] = 5'b00000; w[111][137] = 5'b01111; w[111][138] = 5'b01111; w[111][139] = 5'b01111; w[111][140] = 5'b01111; w[111][141] = 5'b01111; w[111][142] = 5'b01111; w[111][143] = 5'b00000; w[111][144] = 5'b00000; w[111][145] = 5'b01111; w[111][146] = 5'b00000; w[111][147] = 5'b10000; w[111][148] = 5'b01111; w[111][149] = 5'b00000; w[111][150] = 5'b00000; w[111][151] = 5'b01111; w[111][152] = 5'b01111; w[111][153] = 5'b01111; w[111][154] = 5'b01111; w[111][155] = 5'b01111; w[111][156] = 5'b01111; w[111][157] = 5'b00000; w[111][158] = 5'b00000; w[111][159] = 5'b00000; w[111][160] = 5'b10000; w[111][161] = 5'b10000; w[111][162] = 5'b10000; w[111][163] = 5'b00000; w[111][164] = 5'b00000; w[111][165] = 5'b01111; w[111][166] = 5'b01111; w[111][167] = 5'b01111; w[111][168] = 5'b01111; w[111][169] = 5'b01111; w[111][170] = 5'b01111; w[111][171] = 5'b01111; w[111][172] = 5'b00000; w[111][173] = 5'b00000; w[111][174] = 5'b10000; w[111][175] = 5'b10000; w[111][176] = 5'b10000; w[111][177] = 5'b00000; w[111][178] = 5'b01111; w[111][179] = 5'b01111; w[111][180] = 5'b01111; w[111][181] = 5'b01111; w[111][182] = 5'b01111; w[111][183] = 5'b01111; w[111][184] = 5'b01111; w[111][185] = 5'b01111; w[111][186] = 5'b01111; w[111][187] = 5'b01111; w[111][188] = 5'b01111; w[111][189] = 5'b01111; w[111][190] = 5'b01111; w[111][191] = 5'b01111; w[111][192] = 5'b01111; w[111][193] = 5'b01111; w[111][194] = 5'b01111; w[111][195] = 5'b01111; w[111][196] = 5'b01111; w[111][197] = 5'b01111; w[111][198] = 5'b01111; w[111][199] = 5'b01111; w[111][200] = 5'b01111; w[111][201] = 5'b01111; w[111][202] = 5'b01111; w[111][203] = 5'b01111; w[111][204] = 5'b01111; w[111][205] = 5'b01111; w[111][206] = 5'b01111; w[111][207] = 5'b01111; w[111][208] = 5'b01111; w[111][209] = 5'b01111; 
w[112][0] = 5'b01111; w[112][1] = 5'b01111; w[112][2] = 5'b01111; w[112][3] = 5'b01111; w[112][4] = 5'b01111; w[112][5] = 5'b01111; w[112][6] = 5'b01111; w[112][7] = 5'b01111; w[112][8] = 5'b01111; w[112][9] = 5'b01111; w[112][10] = 5'b01111; w[112][11] = 5'b01111; w[112][12] = 5'b01111; w[112][13] = 5'b01111; w[112][14] = 5'b01111; w[112][15] = 5'b01111; w[112][16] = 5'b01111; w[112][17] = 5'b01111; w[112][18] = 5'b01111; w[112][19] = 5'b01111; w[112][20] = 5'b01111; w[112][21] = 5'b01111; w[112][22] = 5'b01111; w[112][23] = 5'b01111; w[112][24] = 5'b01111; w[112][25] = 5'b01111; w[112][26] = 5'b01111; w[112][27] = 5'b01111; w[112][28] = 5'b01111; w[112][29] = 5'b01111; w[112][30] = 5'b01111; w[112][31] = 5'b00000; w[112][32] = 5'b10000; w[112][33] = 5'b10000; w[112][34] = 5'b10000; w[112][35] = 5'b10000; w[112][36] = 5'b10000; w[112][37] = 5'b10000; w[112][38] = 5'b00000; w[112][39] = 5'b01111; w[112][40] = 5'b01111; w[112][41] = 5'b01111; w[112][42] = 5'b01111; w[112][43] = 5'b01111; w[112][44] = 5'b01111; w[112][45] = 5'b10000; w[112][46] = 5'b10000; w[112][47] = 5'b10000; w[112][48] = 5'b10000; w[112][49] = 5'b10000; w[112][50] = 5'b10000; w[112][51] = 5'b10000; w[112][52] = 5'b10000; w[112][53] = 5'b01111; w[112][54] = 5'b01111; w[112][55] = 5'b01111; w[112][56] = 5'b01111; w[112][57] = 5'b01111; w[112][58] = 5'b01111; w[112][59] = 5'b00000; w[112][60] = 5'b00000; w[112][61] = 5'b01111; w[112][62] = 5'b10000; w[112][63] = 5'b00000; w[112][64] = 5'b01111; w[112][65] = 5'b00000; w[112][66] = 5'b00000; w[112][67] = 5'b01111; w[112][68] = 5'b01111; w[112][69] = 5'b01111; w[112][70] = 5'b01111; w[112][71] = 5'b01111; w[112][72] = 5'b01111; w[112][73] = 5'b00000; w[112][74] = 5'b01111; w[112][75] = 5'b01111; w[112][76] = 5'b10000; w[112][77] = 5'b00000; w[112][78] = 5'b01111; w[112][79] = 5'b01111; w[112][80] = 5'b00000; w[112][81] = 5'b01111; w[112][82] = 5'b01111; w[112][83] = 5'b01111; w[112][84] = 5'b01111; w[112][85] = 5'b01111; w[112][86] = 5'b01111; w[112][87] = 5'b00000; w[112][88] = 5'b01111; w[112][89] = 5'b01111; w[112][90] = 5'b10000; w[112][91] = 5'b10000; w[112][92] = 5'b01111; w[112][93] = 5'b01111; w[112][94] = 5'b01111; w[112][95] = 5'b01111; w[112][96] = 5'b01111; w[112][97] = 5'b01111; w[112][98] = 5'b01111; w[112][99] = 5'b01111; w[112][100] = 5'b01111; w[112][101] = 5'b00000; w[112][102] = 5'b01111; w[112][103] = 5'b01111; w[112][104] = 5'b10000; w[112][105] = 5'b10000; w[112][106] = 5'b01111; w[112][107] = 5'b00000; w[112][108] = 5'b00000; w[112][109] = 5'b01111; w[112][110] = 5'b01111; w[112][111] = 5'b01111; w[112][112] = 5'b00000; w[112][113] = 5'b01111; w[112][114] = 5'b01111; w[112][115] = 5'b00000; w[112][116] = 5'b01111; w[112][117] = 5'b01111; w[112][118] = 5'b10000; w[112][119] = 5'b10000; w[112][120] = 5'b00000; w[112][121] = 5'b00000; w[112][122] = 5'b00000; w[112][123] = 5'b01111; w[112][124] = 5'b01111; w[112][125] = 5'b01111; w[112][126] = 5'b01111; w[112][127] = 5'b01111; w[112][128] = 5'b01111; w[112][129] = 5'b00000; w[112][130] = 5'b01111; w[112][131] = 5'b01111; w[112][132] = 5'b00000; w[112][133] = 5'b10000; w[112][134] = 5'b01111; w[112][135] = 5'b01111; w[112][136] = 5'b00000; w[112][137] = 5'b01111; w[112][138] = 5'b01111; w[112][139] = 5'b01111; w[112][140] = 5'b01111; w[112][141] = 5'b01111; w[112][142] = 5'b01111; w[112][143] = 5'b00000; w[112][144] = 5'b00000; w[112][145] = 5'b01111; w[112][146] = 5'b00000; w[112][147] = 5'b10000; w[112][148] = 5'b01111; w[112][149] = 5'b00000; w[112][150] = 5'b00000; w[112][151] = 5'b01111; w[112][152] = 5'b01111; w[112][153] = 5'b01111; w[112][154] = 5'b01111; w[112][155] = 5'b01111; w[112][156] = 5'b01111; w[112][157] = 5'b00000; w[112][158] = 5'b00000; w[112][159] = 5'b00000; w[112][160] = 5'b10000; w[112][161] = 5'b10000; w[112][162] = 5'b10000; w[112][163] = 5'b00000; w[112][164] = 5'b00000; w[112][165] = 5'b01111; w[112][166] = 5'b01111; w[112][167] = 5'b01111; w[112][168] = 5'b01111; w[112][169] = 5'b01111; w[112][170] = 5'b01111; w[112][171] = 5'b01111; w[112][172] = 5'b00000; w[112][173] = 5'b00000; w[112][174] = 5'b10000; w[112][175] = 5'b10000; w[112][176] = 5'b10000; w[112][177] = 5'b00000; w[112][178] = 5'b01111; w[112][179] = 5'b01111; w[112][180] = 5'b01111; w[112][181] = 5'b01111; w[112][182] = 5'b01111; w[112][183] = 5'b01111; w[112][184] = 5'b01111; w[112][185] = 5'b01111; w[112][186] = 5'b01111; w[112][187] = 5'b01111; w[112][188] = 5'b01111; w[112][189] = 5'b01111; w[112][190] = 5'b01111; w[112][191] = 5'b01111; w[112][192] = 5'b01111; w[112][193] = 5'b01111; w[112][194] = 5'b01111; w[112][195] = 5'b01111; w[112][196] = 5'b01111; w[112][197] = 5'b01111; w[112][198] = 5'b01111; w[112][199] = 5'b01111; w[112][200] = 5'b01111; w[112][201] = 5'b01111; w[112][202] = 5'b01111; w[112][203] = 5'b01111; w[112][204] = 5'b01111; w[112][205] = 5'b01111; w[112][206] = 5'b01111; w[112][207] = 5'b01111; w[112][208] = 5'b01111; w[112][209] = 5'b01111; 
w[113][0] = 5'b01111; w[113][1] = 5'b01111; w[113][2] = 5'b01111; w[113][3] = 5'b01111; w[113][4] = 5'b01111; w[113][5] = 5'b01111; w[113][6] = 5'b01111; w[113][7] = 5'b01111; w[113][8] = 5'b01111; w[113][9] = 5'b01111; w[113][10] = 5'b01111; w[113][11] = 5'b01111; w[113][12] = 5'b01111; w[113][13] = 5'b01111; w[113][14] = 5'b01111; w[113][15] = 5'b01111; w[113][16] = 5'b01111; w[113][17] = 5'b01111; w[113][18] = 5'b01111; w[113][19] = 5'b01111; w[113][20] = 5'b01111; w[113][21] = 5'b01111; w[113][22] = 5'b01111; w[113][23] = 5'b01111; w[113][24] = 5'b01111; w[113][25] = 5'b01111; w[113][26] = 5'b01111; w[113][27] = 5'b01111; w[113][28] = 5'b01111; w[113][29] = 5'b01111; w[113][30] = 5'b01111; w[113][31] = 5'b00000; w[113][32] = 5'b10000; w[113][33] = 5'b10000; w[113][34] = 5'b10000; w[113][35] = 5'b10000; w[113][36] = 5'b10000; w[113][37] = 5'b10000; w[113][38] = 5'b00000; w[113][39] = 5'b01111; w[113][40] = 5'b01111; w[113][41] = 5'b01111; w[113][42] = 5'b01111; w[113][43] = 5'b01111; w[113][44] = 5'b01111; w[113][45] = 5'b10000; w[113][46] = 5'b10000; w[113][47] = 5'b10000; w[113][48] = 5'b10000; w[113][49] = 5'b10000; w[113][50] = 5'b10000; w[113][51] = 5'b10000; w[113][52] = 5'b10000; w[113][53] = 5'b01111; w[113][54] = 5'b01111; w[113][55] = 5'b01111; w[113][56] = 5'b01111; w[113][57] = 5'b01111; w[113][58] = 5'b01111; w[113][59] = 5'b00000; w[113][60] = 5'b00000; w[113][61] = 5'b01111; w[113][62] = 5'b10000; w[113][63] = 5'b00000; w[113][64] = 5'b01111; w[113][65] = 5'b00000; w[113][66] = 5'b00000; w[113][67] = 5'b01111; w[113][68] = 5'b01111; w[113][69] = 5'b01111; w[113][70] = 5'b01111; w[113][71] = 5'b01111; w[113][72] = 5'b01111; w[113][73] = 5'b00000; w[113][74] = 5'b01111; w[113][75] = 5'b01111; w[113][76] = 5'b10000; w[113][77] = 5'b00000; w[113][78] = 5'b01111; w[113][79] = 5'b01111; w[113][80] = 5'b00000; w[113][81] = 5'b01111; w[113][82] = 5'b01111; w[113][83] = 5'b01111; w[113][84] = 5'b01111; w[113][85] = 5'b01111; w[113][86] = 5'b01111; w[113][87] = 5'b00000; w[113][88] = 5'b01111; w[113][89] = 5'b01111; w[113][90] = 5'b10000; w[113][91] = 5'b10000; w[113][92] = 5'b01111; w[113][93] = 5'b01111; w[113][94] = 5'b01111; w[113][95] = 5'b01111; w[113][96] = 5'b01111; w[113][97] = 5'b01111; w[113][98] = 5'b01111; w[113][99] = 5'b01111; w[113][100] = 5'b01111; w[113][101] = 5'b00000; w[113][102] = 5'b01111; w[113][103] = 5'b01111; w[113][104] = 5'b10000; w[113][105] = 5'b10000; w[113][106] = 5'b01111; w[113][107] = 5'b00000; w[113][108] = 5'b00000; w[113][109] = 5'b01111; w[113][110] = 5'b01111; w[113][111] = 5'b01111; w[113][112] = 5'b01111; w[113][113] = 5'b00000; w[113][114] = 5'b01111; w[113][115] = 5'b00000; w[113][116] = 5'b01111; w[113][117] = 5'b01111; w[113][118] = 5'b10000; w[113][119] = 5'b10000; w[113][120] = 5'b00000; w[113][121] = 5'b00000; w[113][122] = 5'b00000; w[113][123] = 5'b01111; w[113][124] = 5'b01111; w[113][125] = 5'b01111; w[113][126] = 5'b01111; w[113][127] = 5'b01111; w[113][128] = 5'b01111; w[113][129] = 5'b00000; w[113][130] = 5'b01111; w[113][131] = 5'b01111; w[113][132] = 5'b00000; w[113][133] = 5'b10000; w[113][134] = 5'b01111; w[113][135] = 5'b01111; w[113][136] = 5'b00000; w[113][137] = 5'b01111; w[113][138] = 5'b01111; w[113][139] = 5'b01111; w[113][140] = 5'b01111; w[113][141] = 5'b01111; w[113][142] = 5'b01111; w[113][143] = 5'b00000; w[113][144] = 5'b00000; w[113][145] = 5'b01111; w[113][146] = 5'b00000; w[113][147] = 5'b10000; w[113][148] = 5'b01111; w[113][149] = 5'b00000; w[113][150] = 5'b00000; w[113][151] = 5'b01111; w[113][152] = 5'b01111; w[113][153] = 5'b01111; w[113][154] = 5'b01111; w[113][155] = 5'b01111; w[113][156] = 5'b01111; w[113][157] = 5'b00000; w[113][158] = 5'b00000; w[113][159] = 5'b00000; w[113][160] = 5'b10000; w[113][161] = 5'b10000; w[113][162] = 5'b10000; w[113][163] = 5'b00000; w[113][164] = 5'b00000; w[113][165] = 5'b01111; w[113][166] = 5'b01111; w[113][167] = 5'b01111; w[113][168] = 5'b01111; w[113][169] = 5'b01111; w[113][170] = 5'b01111; w[113][171] = 5'b01111; w[113][172] = 5'b00000; w[113][173] = 5'b00000; w[113][174] = 5'b10000; w[113][175] = 5'b10000; w[113][176] = 5'b10000; w[113][177] = 5'b00000; w[113][178] = 5'b01111; w[113][179] = 5'b01111; w[113][180] = 5'b01111; w[113][181] = 5'b01111; w[113][182] = 5'b01111; w[113][183] = 5'b01111; w[113][184] = 5'b01111; w[113][185] = 5'b01111; w[113][186] = 5'b01111; w[113][187] = 5'b01111; w[113][188] = 5'b01111; w[113][189] = 5'b01111; w[113][190] = 5'b01111; w[113][191] = 5'b01111; w[113][192] = 5'b01111; w[113][193] = 5'b01111; w[113][194] = 5'b01111; w[113][195] = 5'b01111; w[113][196] = 5'b01111; w[113][197] = 5'b01111; w[113][198] = 5'b01111; w[113][199] = 5'b01111; w[113][200] = 5'b01111; w[113][201] = 5'b01111; w[113][202] = 5'b01111; w[113][203] = 5'b01111; w[113][204] = 5'b01111; w[113][205] = 5'b01111; w[113][206] = 5'b01111; w[113][207] = 5'b01111; w[113][208] = 5'b01111; w[113][209] = 5'b01111; 
w[114][0] = 5'b01111; w[114][1] = 5'b01111; w[114][2] = 5'b01111; w[114][3] = 5'b01111; w[114][4] = 5'b01111; w[114][5] = 5'b01111; w[114][6] = 5'b01111; w[114][7] = 5'b01111; w[114][8] = 5'b01111; w[114][9] = 5'b01111; w[114][10] = 5'b01111; w[114][11] = 5'b01111; w[114][12] = 5'b01111; w[114][13] = 5'b01111; w[114][14] = 5'b01111; w[114][15] = 5'b01111; w[114][16] = 5'b01111; w[114][17] = 5'b01111; w[114][18] = 5'b01111; w[114][19] = 5'b01111; w[114][20] = 5'b01111; w[114][21] = 5'b01111; w[114][22] = 5'b01111; w[114][23] = 5'b01111; w[114][24] = 5'b01111; w[114][25] = 5'b01111; w[114][26] = 5'b01111; w[114][27] = 5'b01111; w[114][28] = 5'b01111; w[114][29] = 5'b01111; w[114][30] = 5'b00000; w[114][31] = 5'b10000; w[114][32] = 5'b00000; w[114][33] = 5'b10000; w[114][34] = 5'b00000; w[114][35] = 5'b00000; w[114][36] = 5'b00000; w[114][37] = 5'b00000; w[114][38] = 5'b10000; w[114][39] = 5'b00000; w[114][40] = 5'b01111; w[114][41] = 5'b01111; w[114][42] = 5'b01111; w[114][43] = 5'b01111; w[114][44] = 5'b00000; w[114][45] = 5'b00000; w[114][46] = 5'b00000; w[114][47] = 5'b10000; w[114][48] = 5'b00000; w[114][49] = 5'b00000; w[114][50] = 5'b00000; w[114][51] = 5'b00000; w[114][52] = 5'b00000; w[114][53] = 5'b00000; w[114][54] = 5'b01111; w[114][55] = 5'b01111; w[114][56] = 5'b01111; w[114][57] = 5'b01111; w[114][58] = 5'b01111; w[114][59] = 5'b01111; w[114][60] = 5'b01111; w[114][61] = 5'b00000; w[114][62] = 5'b10000; w[114][63] = 5'b10000; w[114][64] = 5'b01111; w[114][65] = 5'b01111; w[114][66] = 5'b01111; w[114][67] = 5'b01111; w[114][68] = 5'b01111; w[114][69] = 5'b01111; w[114][70] = 5'b01111; w[114][71] = 5'b01111; w[114][72] = 5'b01111; w[114][73] = 5'b01111; w[114][74] = 5'b00000; w[114][75] = 5'b00000; w[114][76] = 5'b10000; w[114][77] = 5'b10000; w[114][78] = 5'b01111; w[114][79] = 5'b00000; w[114][80] = 5'b01111; w[114][81] = 5'b01111; w[114][82] = 5'b01111; w[114][83] = 5'b01111; w[114][84] = 5'b01111; w[114][85] = 5'b01111; w[114][86] = 5'b01111; w[114][87] = 5'b01111; w[114][88] = 5'b00000; w[114][89] = 5'b00000; w[114][90] = 5'b10000; w[114][91] = 5'b10000; w[114][92] = 5'b01111; w[114][93] = 5'b00000; w[114][94] = 5'b00000; w[114][95] = 5'b01111; w[114][96] = 5'b01111; w[114][97] = 5'b01111; w[114][98] = 5'b01111; w[114][99] = 5'b01111; w[114][100] = 5'b01111; w[114][101] = 5'b01111; w[114][102] = 5'b00000; w[114][103] = 5'b01111; w[114][104] = 5'b10000; w[114][105] = 5'b10000; w[114][106] = 5'b01111; w[114][107] = 5'b01111; w[114][108] = 5'b01111; w[114][109] = 5'b01111; w[114][110] = 5'b01111; w[114][111] = 5'b01111; w[114][112] = 5'b01111; w[114][113] = 5'b01111; w[114][114] = 5'b00000; w[114][115] = 5'b01111; w[114][116] = 5'b00000; w[114][117] = 5'b01111; w[114][118] = 5'b10000; w[114][119] = 5'b10000; w[114][120] = 5'b01111; w[114][121] = 5'b01111; w[114][122] = 5'b01111; w[114][123] = 5'b01111; w[114][124] = 5'b01111; w[114][125] = 5'b01111; w[114][126] = 5'b01111; w[114][127] = 5'b01111; w[114][128] = 5'b01111; w[114][129] = 5'b01111; w[114][130] = 5'b00000; w[114][131] = 5'b01111; w[114][132] = 5'b10000; w[114][133] = 5'b10000; w[114][134] = 5'b00000; w[114][135] = 5'b00000; w[114][136] = 5'b01111; w[114][137] = 5'b01111; w[114][138] = 5'b01111; w[114][139] = 5'b01111; w[114][140] = 5'b01111; w[114][141] = 5'b01111; w[114][142] = 5'b01111; w[114][143] = 5'b01111; w[114][144] = 5'b01111; w[114][145] = 5'b01111; w[114][146] = 5'b10000; w[114][147] = 5'b10000; w[114][148] = 5'b00000; w[114][149] = 5'b01111; w[114][150] = 5'b01111; w[114][151] = 5'b01111; w[114][152] = 5'b01111; w[114][153] = 5'b01111; w[114][154] = 5'b01111; w[114][155] = 5'b01111; w[114][156] = 5'b01111; w[114][157] = 5'b01111; w[114][158] = 5'b01111; w[114][159] = 5'b01111; w[114][160] = 5'b00000; w[114][161] = 5'b00000; w[114][162] = 5'b00000; w[114][163] = 5'b01111; w[114][164] = 5'b01111; w[114][165] = 5'b01111; w[114][166] = 5'b01111; w[114][167] = 5'b01111; w[114][168] = 5'b01111; w[114][169] = 5'b01111; w[114][170] = 5'b01111; w[114][171] = 5'b00000; w[114][172] = 5'b01111; w[114][173] = 5'b01111; w[114][174] = 5'b00000; w[114][175] = 5'b00000; w[114][176] = 5'b00000; w[114][177] = 5'b01111; w[114][178] = 5'b00000; w[114][179] = 5'b01111; w[114][180] = 5'b01111; w[114][181] = 5'b01111; w[114][182] = 5'b01111; w[114][183] = 5'b01111; w[114][184] = 5'b01111; w[114][185] = 5'b01111; w[114][186] = 5'b01111; w[114][187] = 5'b01111; w[114][188] = 5'b01111; w[114][189] = 5'b01111; w[114][190] = 5'b01111; w[114][191] = 5'b01111; w[114][192] = 5'b01111; w[114][193] = 5'b01111; w[114][194] = 5'b01111; w[114][195] = 5'b01111; w[114][196] = 5'b01111; w[114][197] = 5'b01111; w[114][198] = 5'b01111; w[114][199] = 5'b01111; w[114][200] = 5'b01111; w[114][201] = 5'b01111; w[114][202] = 5'b01111; w[114][203] = 5'b01111; w[114][204] = 5'b01111; w[114][205] = 5'b01111; w[114][206] = 5'b01111; w[114][207] = 5'b01111; w[114][208] = 5'b01111; w[114][209] = 5'b01111; 
w[115][0] = 5'b00000; w[115][1] = 5'b00000; w[115][2] = 5'b00000; w[115][3] = 5'b00000; w[115][4] = 5'b00000; w[115][5] = 5'b00000; w[115][6] = 5'b00000; w[115][7] = 5'b00000; w[115][8] = 5'b00000; w[115][9] = 5'b00000; w[115][10] = 5'b00000; w[115][11] = 5'b00000; w[115][12] = 5'b00000; w[115][13] = 5'b00000; w[115][14] = 5'b00000; w[115][15] = 5'b00000; w[115][16] = 5'b00000; w[115][17] = 5'b00000; w[115][18] = 5'b00000; w[115][19] = 5'b00000; w[115][20] = 5'b00000; w[115][21] = 5'b00000; w[115][22] = 5'b00000; w[115][23] = 5'b00000; w[115][24] = 5'b00000; w[115][25] = 5'b00000; w[115][26] = 5'b00000; w[115][27] = 5'b00000; w[115][28] = 5'b00000; w[115][29] = 5'b00000; w[115][30] = 5'b10000; w[115][31] = 5'b00000; w[115][32] = 5'b01111; w[115][33] = 5'b00000; w[115][34] = 5'b10000; w[115][35] = 5'b10000; w[115][36] = 5'b10000; w[115][37] = 5'b01111; w[115][38] = 5'b00000; w[115][39] = 5'b10000; w[115][40] = 5'b00000; w[115][41] = 5'b00000; w[115][42] = 5'b00000; w[115][43] = 5'b00000; w[115][44] = 5'b10000; w[115][45] = 5'b01111; w[115][46] = 5'b01111; w[115][47] = 5'b00000; w[115][48] = 5'b10000; w[115][49] = 5'b10000; w[115][50] = 5'b10000; w[115][51] = 5'b01111; w[115][52] = 5'b01111; w[115][53] = 5'b10000; w[115][54] = 5'b00000; w[115][55] = 5'b00000; w[115][56] = 5'b00000; w[115][57] = 5'b00000; w[115][58] = 5'b01111; w[115][59] = 5'b01111; w[115][60] = 5'b01111; w[115][61] = 5'b01111; w[115][62] = 5'b10000; w[115][63] = 5'b10000; w[115][64] = 5'b00000; w[115][65] = 5'b01111; w[115][66] = 5'b01111; w[115][67] = 5'b01111; w[115][68] = 5'b00000; w[115][69] = 5'b00000; w[115][70] = 5'b00000; w[115][71] = 5'b00000; w[115][72] = 5'b01111; w[115][73] = 5'b01111; w[115][74] = 5'b01111; w[115][75] = 5'b01111; w[115][76] = 5'b10000; w[115][77] = 5'b10000; w[115][78] = 5'b00000; w[115][79] = 5'b01111; w[115][80] = 5'b01111; w[115][81] = 5'b01111; w[115][82] = 5'b00000; w[115][83] = 5'b00000; w[115][84] = 5'b00000; w[115][85] = 5'b00000; w[115][86] = 5'b01111; w[115][87] = 5'b01111; w[115][88] = 5'b01111; w[115][89] = 5'b01111; w[115][90] = 5'b10000; w[115][91] = 5'b10000; w[115][92] = 5'b00000; w[115][93] = 5'b01111; w[115][94] = 5'b01111; w[115][95] = 5'b00000; w[115][96] = 5'b00000; w[115][97] = 5'b00000; w[115][98] = 5'b00000; w[115][99] = 5'b00000; w[115][100] = 5'b01111; w[115][101] = 5'b01111; w[115][102] = 5'b01111; w[115][103] = 5'b00000; w[115][104] = 5'b10000; w[115][105] = 5'b10000; w[115][106] = 5'b01111; w[115][107] = 5'b01111; w[115][108] = 5'b01111; w[115][109] = 5'b01111; w[115][110] = 5'b00000; w[115][111] = 5'b00000; w[115][112] = 5'b00000; w[115][113] = 5'b00000; w[115][114] = 5'b01111; w[115][115] = 5'b00000; w[115][116] = 5'b01111; w[115][117] = 5'b00000; w[115][118] = 5'b10000; w[115][119] = 5'b10000; w[115][120] = 5'b01111; w[115][121] = 5'b01111; w[115][122] = 5'b01111; w[115][123] = 5'b01111; w[115][124] = 5'b00000; w[115][125] = 5'b00000; w[115][126] = 5'b00000; w[115][127] = 5'b00000; w[115][128] = 5'b01111; w[115][129] = 5'b01111; w[115][130] = 5'b01111; w[115][131] = 5'b00000; w[115][132] = 5'b10000; w[115][133] = 5'b10000; w[115][134] = 5'b01111; w[115][135] = 5'b01111; w[115][136] = 5'b01111; w[115][137] = 5'b01111; w[115][138] = 5'b00000; w[115][139] = 5'b00000; w[115][140] = 5'b00000; w[115][141] = 5'b00000; w[115][142] = 5'b01111; w[115][143] = 5'b01111; w[115][144] = 5'b01111; w[115][145] = 5'b00000; w[115][146] = 5'b10000; w[115][147] = 5'b10000; w[115][148] = 5'b01111; w[115][149] = 5'b01111; w[115][150] = 5'b01111; w[115][151] = 5'b01111; w[115][152] = 5'b00000; w[115][153] = 5'b00000; w[115][154] = 5'b00000; w[115][155] = 5'b00000; w[115][156] = 5'b00000; w[115][157] = 5'b01111; w[115][158] = 5'b01111; w[115][159] = 5'b00000; w[115][160] = 5'b10000; w[115][161] = 5'b10000; w[115][162] = 5'b01111; w[115][163] = 5'b01111; w[115][164] = 5'b01111; w[115][165] = 5'b00000; w[115][166] = 5'b00000; w[115][167] = 5'b00000; w[115][168] = 5'b00000; w[115][169] = 5'b00000; w[115][170] = 5'b00000; w[115][171] = 5'b01111; w[115][172] = 5'b01111; w[115][173] = 5'b00000; w[115][174] = 5'b10000; w[115][175] = 5'b10000; w[115][176] = 5'b01111; w[115][177] = 5'b01111; w[115][178] = 5'b01111; w[115][179] = 5'b00000; w[115][180] = 5'b00000; w[115][181] = 5'b00000; w[115][182] = 5'b00000; w[115][183] = 5'b00000; w[115][184] = 5'b00000; w[115][185] = 5'b00000; w[115][186] = 5'b00000; w[115][187] = 5'b00000; w[115][188] = 5'b00000; w[115][189] = 5'b00000; w[115][190] = 5'b00000; w[115][191] = 5'b00000; w[115][192] = 5'b00000; w[115][193] = 5'b00000; w[115][194] = 5'b00000; w[115][195] = 5'b00000; w[115][196] = 5'b00000; w[115][197] = 5'b00000; w[115][198] = 5'b00000; w[115][199] = 5'b00000; w[115][200] = 5'b00000; w[115][201] = 5'b00000; w[115][202] = 5'b00000; w[115][203] = 5'b00000; w[115][204] = 5'b00000; w[115][205] = 5'b00000; w[115][206] = 5'b00000; w[115][207] = 5'b00000; w[115][208] = 5'b00000; w[115][209] = 5'b00000; 
w[116][0] = 5'b01111; w[116][1] = 5'b01111; w[116][2] = 5'b01111; w[116][3] = 5'b01111; w[116][4] = 5'b01111; w[116][5] = 5'b01111; w[116][6] = 5'b01111; w[116][7] = 5'b01111; w[116][8] = 5'b01111; w[116][9] = 5'b01111; w[116][10] = 5'b01111; w[116][11] = 5'b01111; w[116][12] = 5'b01111; w[116][13] = 5'b01111; w[116][14] = 5'b01111; w[116][15] = 5'b01111; w[116][16] = 5'b01111; w[116][17] = 5'b01111; w[116][18] = 5'b01111; w[116][19] = 5'b01111; w[116][20] = 5'b01111; w[116][21] = 5'b01111; w[116][22] = 5'b01111; w[116][23] = 5'b01111; w[116][24] = 5'b01111; w[116][25] = 5'b01111; w[116][26] = 5'b01111; w[116][27] = 5'b01111; w[116][28] = 5'b01111; w[116][29] = 5'b01111; w[116][30] = 5'b00000; w[116][31] = 5'b01111; w[116][32] = 5'b00000; w[116][33] = 5'b10000; w[116][34] = 5'b10000; w[116][35] = 5'b10000; w[116][36] = 5'b10000; w[116][37] = 5'b00000; w[116][38] = 5'b01111; w[116][39] = 5'b00000; w[116][40] = 5'b01111; w[116][41] = 5'b01111; w[116][42] = 5'b01111; w[116][43] = 5'b01111; w[116][44] = 5'b00000; w[116][45] = 5'b00000; w[116][46] = 5'b00000; w[116][47] = 5'b10000; w[116][48] = 5'b10000; w[116][49] = 5'b10000; w[116][50] = 5'b10000; w[116][51] = 5'b00000; w[116][52] = 5'b00000; w[116][53] = 5'b00000; w[116][54] = 5'b01111; w[116][55] = 5'b01111; w[116][56] = 5'b01111; w[116][57] = 5'b01111; w[116][58] = 5'b00000; w[116][59] = 5'b01111; w[116][60] = 5'b01111; w[116][61] = 5'b01111; w[116][62] = 5'b00000; w[116][63] = 5'b10000; w[116][64] = 5'b01111; w[116][65] = 5'b01111; w[116][66] = 5'b01111; w[116][67] = 5'b00000; w[116][68] = 5'b01111; w[116][69] = 5'b01111; w[116][70] = 5'b01111; w[116][71] = 5'b01111; w[116][72] = 5'b00000; w[116][73] = 5'b01111; w[116][74] = 5'b01111; w[116][75] = 5'b01111; w[116][76] = 5'b00000; w[116][77] = 5'b10000; w[116][78] = 5'b01111; w[116][79] = 5'b01111; w[116][80] = 5'b01111; w[116][81] = 5'b00000; w[116][82] = 5'b01111; w[116][83] = 5'b01111; w[116][84] = 5'b01111; w[116][85] = 5'b01111; w[116][86] = 5'b00000; w[116][87] = 5'b01111; w[116][88] = 5'b01111; w[116][89] = 5'b01111; w[116][90] = 5'b00000; w[116][91] = 5'b00000; w[116][92] = 5'b01111; w[116][93] = 5'b01111; w[116][94] = 5'b01111; w[116][95] = 5'b01111; w[116][96] = 5'b01111; w[116][97] = 5'b01111; w[116][98] = 5'b01111; w[116][99] = 5'b01111; w[116][100] = 5'b00000; w[116][101] = 5'b01111; w[116][102] = 5'b01111; w[116][103] = 5'b01111; w[116][104] = 5'b00000; w[116][105] = 5'b00000; w[116][106] = 5'b00000; w[116][107] = 5'b01111; w[116][108] = 5'b01111; w[116][109] = 5'b00000; w[116][110] = 5'b01111; w[116][111] = 5'b01111; w[116][112] = 5'b01111; w[116][113] = 5'b01111; w[116][114] = 5'b00000; w[116][115] = 5'b01111; w[116][116] = 5'b00000; w[116][117] = 5'b01111; w[116][118] = 5'b00000; w[116][119] = 5'b00000; w[116][120] = 5'b01111; w[116][121] = 5'b01111; w[116][122] = 5'b01111; w[116][123] = 5'b00000; w[116][124] = 5'b01111; w[116][125] = 5'b01111; w[116][126] = 5'b01111; w[116][127] = 5'b01111; w[116][128] = 5'b00000; w[116][129] = 5'b01111; w[116][130] = 5'b01111; w[116][131] = 5'b01111; w[116][132] = 5'b10000; w[116][133] = 5'b00000; w[116][134] = 5'b01111; w[116][135] = 5'b01111; w[116][136] = 5'b01111; w[116][137] = 5'b00000; w[116][138] = 5'b01111; w[116][139] = 5'b01111; w[116][140] = 5'b01111; w[116][141] = 5'b01111; w[116][142] = 5'b00000; w[116][143] = 5'b01111; w[116][144] = 5'b01111; w[116][145] = 5'b01111; w[116][146] = 5'b10000; w[116][147] = 5'b00000; w[116][148] = 5'b01111; w[116][149] = 5'b01111; w[116][150] = 5'b01111; w[116][151] = 5'b00000; w[116][152] = 5'b01111; w[116][153] = 5'b01111; w[116][154] = 5'b01111; w[116][155] = 5'b01111; w[116][156] = 5'b01111; w[116][157] = 5'b01111; w[116][158] = 5'b01111; w[116][159] = 5'b10000; w[116][160] = 5'b10000; w[116][161] = 5'b10000; w[116][162] = 5'b00000; w[116][163] = 5'b01111; w[116][164] = 5'b01111; w[116][165] = 5'b01111; w[116][166] = 5'b01111; w[116][167] = 5'b01111; w[116][168] = 5'b01111; w[116][169] = 5'b01111; w[116][170] = 5'b01111; w[116][171] = 5'b01111; w[116][172] = 5'b01111; w[116][173] = 5'b10000; w[116][174] = 5'b10000; w[116][175] = 5'b10000; w[116][176] = 5'b00000; w[116][177] = 5'b01111; w[116][178] = 5'b01111; w[116][179] = 5'b01111; w[116][180] = 5'b01111; w[116][181] = 5'b01111; w[116][182] = 5'b01111; w[116][183] = 5'b01111; w[116][184] = 5'b01111; w[116][185] = 5'b01111; w[116][186] = 5'b01111; w[116][187] = 5'b01111; w[116][188] = 5'b01111; w[116][189] = 5'b01111; w[116][190] = 5'b01111; w[116][191] = 5'b01111; w[116][192] = 5'b01111; w[116][193] = 5'b01111; w[116][194] = 5'b01111; w[116][195] = 5'b01111; w[116][196] = 5'b01111; w[116][197] = 5'b01111; w[116][198] = 5'b01111; w[116][199] = 5'b01111; w[116][200] = 5'b01111; w[116][201] = 5'b01111; w[116][202] = 5'b01111; w[116][203] = 5'b01111; w[116][204] = 5'b01111; w[116][205] = 5'b01111; w[116][206] = 5'b01111; w[116][207] = 5'b01111; w[116][208] = 5'b01111; w[116][209] = 5'b01111; 
w[117][0] = 5'b01111; w[117][1] = 5'b01111; w[117][2] = 5'b01111; w[117][3] = 5'b01111; w[117][4] = 5'b01111; w[117][5] = 5'b01111; w[117][6] = 5'b01111; w[117][7] = 5'b01111; w[117][8] = 5'b01111; w[117][9] = 5'b01111; w[117][10] = 5'b01111; w[117][11] = 5'b01111; w[117][12] = 5'b01111; w[117][13] = 5'b01111; w[117][14] = 5'b01111; w[117][15] = 5'b01111; w[117][16] = 5'b01111; w[117][17] = 5'b01111; w[117][18] = 5'b01111; w[117][19] = 5'b01111; w[117][20] = 5'b01111; w[117][21] = 5'b01111; w[117][22] = 5'b01111; w[117][23] = 5'b01111; w[117][24] = 5'b01111; w[117][25] = 5'b01111; w[117][26] = 5'b01111; w[117][27] = 5'b01111; w[117][28] = 5'b01111; w[117][29] = 5'b01111; w[117][30] = 5'b01111; w[117][31] = 5'b00000; w[117][32] = 5'b10000; w[117][33] = 5'b10000; w[117][34] = 5'b10000; w[117][35] = 5'b10000; w[117][36] = 5'b10000; w[117][37] = 5'b10000; w[117][38] = 5'b00000; w[117][39] = 5'b01111; w[117][40] = 5'b01111; w[117][41] = 5'b01111; w[117][42] = 5'b01111; w[117][43] = 5'b01111; w[117][44] = 5'b01111; w[117][45] = 5'b10000; w[117][46] = 5'b10000; w[117][47] = 5'b10000; w[117][48] = 5'b10000; w[117][49] = 5'b10000; w[117][50] = 5'b10000; w[117][51] = 5'b10000; w[117][52] = 5'b10000; w[117][53] = 5'b01111; w[117][54] = 5'b01111; w[117][55] = 5'b01111; w[117][56] = 5'b01111; w[117][57] = 5'b01111; w[117][58] = 5'b01111; w[117][59] = 5'b00000; w[117][60] = 5'b00000; w[117][61] = 5'b01111; w[117][62] = 5'b10000; w[117][63] = 5'b00000; w[117][64] = 5'b01111; w[117][65] = 5'b00000; w[117][66] = 5'b00000; w[117][67] = 5'b01111; w[117][68] = 5'b01111; w[117][69] = 5'b01111; w[117][70] = 5'b01111; w[117][71] = 5'b01111; w[117][72] = 5'b01111; w[117][73] = 5'b00000; w[117][74] = 5'b01111; w[117][75] = 5'b01111; w[117][76] = 5'b10000; w[117][77] = 5'b00000; w[117][78] = 5'b01111; w[117][79] = 5'b01111; w[117][80] = 5'b00000; w[117][81] = 5'b01111; w[117][82] = 5'b01111; w[117][83] = 5'b01111; w[117][84] = 5'b01111; w[117][85] = 5'b01111; w[117][86] = 5'b01111; w[117][87] = 5'b00000; w[117][88] = 5'b01111; w[117][89] = 5'b01111; w[117][90] = 5'b10000; w[117][91] = 5'b10000; w[117][92] = 5'b01111; w[117][93] = 5'b01111; w[117][94] = 5'b01111; w[117][95] = 5'b01111; w[117][96] = 5'b01111; w[117][97] = 5'b01111; w[117][98] = 5'b01111; w[117][99] = 5'b01111; w[117][100] = 5'b01111; w[117][101] = 5'b00000; w[117][102] = 5'b01111; w[117][103] = 5'b01111; w[117][104] = 5'b10000; w[117][105] = 5'b10000; w[117][106] = 5'b01111; w[117][107] = 5'b00000; w[117][108] = 5'b00000; w[117][109] = 5'b01111; w[117][110] = 5'b01111; w[117][111] = 5'b01111; w[117][112] = 5'b01111; w[117][113] = 5'b01111; w[117][114] = 5'b01111; w[117][115] = 5'b00000; w[117][116] = 5'b01111; w[117][117] = 5'b00000; w[117][118] = 5'b10000; w[117][119] = 5'b10000; w[117][120] = 5'b00000; w[117][121] = 5'b00000; w[117][122] = 5'b00000; w[117][123] = 5'b01111; w[117][124] = 5'b01111; w[117][125] = 5'b01111; w[117][126] = 5'b01111; w[117][127] = 5'b01111; w[117][128] = 5'b01111; w[117][129] = 5'b00000; w[117][130] = 5'b01111; w[117][131] = 5'b01111; w[117][132] = 5'b00000; w[117][133] = 5'b10000; w[117][134] = 5'b01111; w[117][135] = 5'b01111; w[117][136] = 5'b00000; w[117][137] = 5'b01111; w[117][138] = 5'b01111; w[117][139] = 5'b01111; w[117][140] = 5'b01111; w[117][141] = 5'b01111; w[117][142] = 5'b01111; w[117][143] = 5'b00000; w[117][144] = 5'b00000; w[117][145] = 5'b01111; w[117][146] = 5'b00000; w[117][147] = 5'b10000; w[117][148] = 5'b01111; w[117][149] = 5'b00000; w[117][150] = 5'b00000; w[117][151] = 5'b01111; w[117][152] = 5'b01111; w[117][153] = 5'b01111; w[117][154] = 5'b01111; w[117][155] = 5'b01111; w[117][156] = 5'b01111; w[117][157] = 5'b00000; w[117][158] = 5'b00000; w[117][159] = 5'b00000; w[117][160] = 5'b10000; w[117][161] = 5'b10000; w[117][162] = 5'b10000; w[117][163] = 5'b00000; w[117][164] = 5'b00000; w[117][165] = 5'b01111; w[117][166] = 5'b01111; w[117][167] = 5'b01111; w[117][168] = 5'b01111; w[117][169] = 5'b01111; w[117][170] = 5'b01111; w[117][171] = 5'b01111; w[117][172] = 5'b00000; w[117][173] = 5'b00000; w[117][174] = 5'b10000; w[117][175] = 5'b10000; w[117][176] = 5'b10000; w[117][177] = 5'b00000; w[117][178] = 5'b01111; w[117][179] = 5'b01111; w[117][180] = 5'b01111; w[117][181] = 5'b01111; w[117][182] = 5'b01111; w[117][183] = 5'b01111; w[117][184] = 5'b01111; w[117][185] = 5'b01111; w[117][186] = 5'b01111; w[117][187] = 5'b01111; w[117][188] = 5'b01111; w[117][189] = 5'b01111; w[117][190] = 5'b01111; w[117][191] = 5'b01111; w[117][192] = 5'b01111; w[117][193] = 5'b01111; w[117][194] = 5'b01111; w[117][195] = 5'b01111; w[117][196] = 5'b01111; w[117][197] = 5'b01111; w[117][198] = 5'b01111; w[117][199] = 5'b01111; w[117][200] = 5'b01111; w[117][201] = 5'b01111; w[117][202] = 5'b01111; w[117][203] = 5'b01111; w[117][204] = 5'b01111; w[117][205] = 5'b01111; w[117][206] = 5'b01111; w[117][207] = 5'b01111; w[117][208] = 5'b01111; w[117][209] = 5'b01111; 
w[118][0] = 5'b10000; w[118][1] = 5'b10000; w[118][2] = 5'b10000; w[118][3] = 5'b10000; w[118][4] = 5'b10000; w[118][5] = 5'b10000; w[118][6] = 5'b10000; w[118][7] = 5'b10000; w[118][8] = 5'b10000; w[118][9] = 5'b10000; w[118][10] = 5'b10000; w[118][11] = 5'b10000; w[118][12] = 5'b10000; w[118][13] = 5'b10000; w[118][14] = 5'b10000; w[118][15] = 5'b10000; w[118][16] = 5'b10000; w[118][17] = 5'b10000; w[118][18] = 5'b10000; w[118][19] = 5'b10000; w[118][20] = 5'b10000; w[118][21] = 5'b10000; w[118][22] = 5'b10000; w[118][23] = 5'b10000; w[118][24] = 5'b10000; w[118][25] = 5'b10000; w[118][26] = 5'b10000; w[118][27] = 5'b10000; w[118][28] = 5'b10000; w[118][29] = 5'b10000; w[118][30] = 5'b00000; w[118][31] = 5'b01111; w[118][32] = 5'b00000; w[118][33] = 5'b01111; w[118][34] = 5'b00000; w[118][35] = 5'b00000; w[118][36] = 5'b00000; w[118][37] = 5'b00000; w[118][38] = 5'b01111; w[118][39] = 5'b00000; w[118][40] = 5'b10000; w[118][41] = 5'b10000; w[118][42] = 5'b10000; w[118][43] = 5'b10000; w[118][44] = 5'b00000; w[118][45] = 5'b00000; w[118][46] = 5'b00000; w[118][47] = 5'b01111; w[118][48] = 5'b00000; w[118][49] = 5'b00000; w[118][50] = 5'b00000; w[118][51] = 5'b00000; w[118][52] = 5'b00000; w[118][53] = 5'b00000; w[118][54] = 5'b10000; w[118][55] = 5'b10000; w[118][56] = 5'b10000; w[118][57] = 5'b10000; w[118][58] = 5'b10000; w[118][59] = 5'b10000; w[118][60] = 5'b10000; w[118][61] = 5'b00000; w[118][62] = 5'b01111; w[118][63] = 5'b01111; w[118][64] = 5'b10000; w[118][65] = 5'b10000; w[118][66] = 5'b10000; w[118][67] = 5'b10000; w[118][68] = 5'b10000; w[118][69] = 5'b10000; w[118][70] = 5'b10000; w[118][71] = 5'b10000; w[118][72] = 5'b10000; w[118][73] = 5'b10000; w[118][74] = 5'b00000; w[118][75] = 5'b00000; w[118][76] = 5'b01111; w[118][77] = 5'b01111; w[118][78] = 5'b10000; w[118][79] = 5'b00000; w[118][80] = 5'b10000; w[118][81] = 5'b10000; w[118][82] = 5'b10000; w[118][83] = 5'b10000; w[118][84] = 5'b10000; w[118][85] = 5'b10000; w[118][86] = 5'b10000; w[118][87] = 5'b10000; w[118][88] = 5'b00000; w[118][89] = 5'b00000; w[118][90] = 5'b01111; w[118][91] = 5'b01111; w[118][92] = 5'b10000; w[118][93] = 5'b00000; w[118][94] = 5'b00000; w[118][95] = 5'b10000; w[118][96] = 5'b10000; w[118][97] = 5'b10000; w[118][98] = 5'b10000; w[118][99] = 5'b10000; w[118][100] = 5'b10000; w[118][101] = 5'b10000; w[118][102] = 5'b00000; w[118][103] = 5'b10000; w[118][104] = 5'b01111; w[118][105] = 5'b01111; w[118][106] = 5'b10000; w[118][107] = 5'b10000; w[118][108] = 5'b10000; w[118][109] = 5'b10000; w[118][110] = 5'b10000; w[118][111] = 5'b10000; w[118][112] = 5'b10000; w[118][113] = 5'b10000; w[118][114] = 5'b10000; w[118][115] = 5'b10000; w[118][116] = 5'b00000; w[118][117] = 5'b10000; w[118][118] = 5'b00000; w[118][119] = 5'b01111; w[118][120] = 5'b10000; w[118][121] = 5'b10000; w[118][122] = 5'b10000; w[118][123] = 5'b10000; w[118][124] = 5'b10000; w[118][125] = 5'b10000; w[118][126] = 5'b10000; w[118][127] = 5'b10000; w[118][128] = 5'b10000; w[118][129] = 5'b10000; w[118][130] = 5'b00000; w[118][131] = 5'b10000; w[118][132] = 5'b01111; w[118][133] = 5'b01111; w[118][134] = 5'b00000; w[118][135] = 5'b00000; w[118][136] = 5'b10000; w[118][137] = 5'b10000; w[118][138] = 5'b10000; w[118][139] = 5'b10000; w[118][140] = 5'b10000; w[118][141] = 5'b10000; w[118][142] = 5'b10000; w[118][143] = 5'b10000; w[118][144] = 5'b10000; w[118][145] = 5'b10000; w[118][146] = 5'b01111; w[118][147] = 5'b01111; w[118][148] = 5'b00000; w[118][149] = 5'b10000; w[118][150] = 5'b10000; w[118][151] = 5'b10000; w[118][152] = 5'b10000; w[118][153] = 5'b10000; w[118][154] = 5'b10000; w[118][155] = 5'b10000; w[118][156] = 5'b10000; w[118][157] = 5'b10000; w[118][158] = 5'b10000; w[118][159] = 5'b10000; w[118][160] = 5'b00000; w[118][161] = 5'b00000; w[118][162] = 5'b00000; w[118][163] = 5'b10000; w[118][164] = 5'b10000; w[118][165] = 5'b10000; w[118][166] = 5'b10000; w[118][167] = 5'b10000; w[118][168] = 5'b10000; w[118][169] = 5'b10000; w[118][170] = 5'b10000; w[118][171] = 5'b00000; w[118][172] = 5'b10000; w[118][173] = 5'b10000; w[118][174] = 5'b00000; w[118][175] = 5'b00000; w[118][176] = 5'b00000; w[118][177] = 5'b10000; w[118][178] = 5'b00000; w[118][179] = 5'b10000; w[118][180] = 5'b10000; w[118][181] = 5'b10000; w[118][182] = 5'b10000; w[118][183] = 5'b10000; w[118][184] = 5'b10000; w[118][185] = 5'b10000; w[118][186] = 5'b10000; w[118][187] = 5'b10000; w[118][188] = 5'b10000; w[118][189] = 5'b10000; w[118][190] = 5'b10000; w[118][191] = 5'b10000; w[118][192] = 5'b10000; w[118][193] = 5'b10000; w[118][194] = 5'b10000; w[118][195] = 5'b10000; w[118][196] = 5'b10000; w[118][197] = 5'b10000; w[118][198] = 5'b10000; w[118][199] = 5'b10000; w[118][200] = 5'b10000; w[118][201] = 5'b10000; w[118][202] = 5'b10000; w[118][203] = 5'b10000; w[118][204] = 5'b10000; w[118][205] = 5'b10000; w[118][206] = 5'b10000; w[118][207] = 5'b10000; w[118][208] = 5'b10000; w[118][209] = 5'b10000; 
w[119][0] = 5'b10000; w[119][1] = 5'b10000; w[119][2] = 5'b10000; w[119][3] = 5'b10000; w[119][4] = 5'b10000; w[119][5] = 5'b10000; w[119][6] = 5'b10000; w[119][7] = 5'b10000; w[119][8] = 5'b10000; w[119][9] = 5'b10000; w[119][10] = 5'b10000; w[119][11] = 5'b10000; w[119][12] = 5'b10000; w[119][13] = 5'b10000; w[119][14] = 5'b10000; w[119][15] = 5'b10000; w[119][16] = 5'b10000; w[119][17] = 5'b10000; w[119][18] = 5'b10000; w[119][19] = 5'b10000; w[119][20] = 5'b10000; w[119][21] = 5'b10000; w[119][22] = 5'b10000; w[119][23] = 5'b10000; w[119][24] = 5'b10000; w[119][25] = 5'b10000; w[119][26] = 5'b10000; w[119][27] = 5'b10000; w[119][28] = 5'b10000; w[119][29] = 5'b10000; w[119][30] = 5'b00000; w[119][31] = 5'b01111; w[119][32] = 5'b00000; w[119][33] = 5'b01111; w[119][34] = 5'b00000; w[119][35] = 5'b00000; w[119][36] = 5'b00000; w[119][37] = 5'b00000; w[119][38] = 5'b01111; w[119][39] = 5'b00000; w[119][40] = 5'b10000; w[119][41] = 5'b10000; w[119][42] = 5'b10000; w[119][43] = 5'b10000; w[119][44] = 5'b00000; w[119][45] = 5'b00000; w[119][46] = 5'b00000; w[119][47] = 5'b01111; w[119][48] = 5'b00000; w[119][49] = 5'b00000; w[119][50] = 5'b00000; w[119][51] = 5'b00000; w[119][52] = 5'b00000; w[119][53] = 5'b00000; w[119][54] = 5'b10000; w[119][55] = 5'b10000; w[119][56] = 5'b10000; w[119][57] = 5'b10000; w[119][58] = 5'b10000; w[119][59] = 5'b10000; w[119][60] = 5'b10000; w[119][61] = 5'b00000; w[119][62] = 5'b01111; w[119][63] = 5'b01111; w[119][64] = 5'b10000; w[119][65] = 5'b10000; w[119][66] = 5'b10000; w[119][67] = 5'b10000; w[119][68] = 5'b10000; w[119][69] = 5'b10000; w[119][70] = 5'b10000; w[119][71] = 5'b10000; w[119][72] = 5'b10000; w[119][73] = 5'b10000; w[119][74] = 5'b00000; w[119][75] = 5'b00000; w[119][76] = 5'b01111; w[119][77] = 5'b01111; w[119][78] = 5'b10000; w[119][79] = 5'b00000; w[119][80] = 5'b10000; w[119][81] = 5'b10000; w[119][82] = 5'b10000; w[119][83] = 5'b10000; w[119][84] = 5'b10000; w[119][85] = 5'b10000; w[119][86] = 5'b10000; w[119][87] = 5'b10000; w[119][88] = 5'b00000; w[119][89] = 5'b00000; w[119][90] = 5'b01111; w[119][91] = 5'b01111; w[119][92] = 5'b10000; w[119][93] = 5'b00000; w[119][94] = 5'b00000; w[119][95] = 5'b10000; w[119][96] = 5'b10000; w[119][97] = 5'b10000; w[119][98] = 5'b10000; w[119][99] = 5'b10000; w[119][100] = 5'b10000; w[119][101] = 5'b10000; w[119][102] = 5'b00000; w[119][103] = 5'b10000; w[119][104] = 5'b01111; w[119][105] = 5'b01111; w[119][106] = 5'b10000; w[119][107] = 5'b10000; w[119][108] = 5'b10000; w[119][109] = 5'b10000; w[119][110] = 5'b10000; w[119][111] = 5'b10000; w[119][112] = 5'b10000; w[119][113] = 5'b10000; w[119][114] = 5'b10000; w[119][115] = 5'b10000; w[119][116] = 5'b00000; w[119][117] = 5'b10000; w[119][118] = 5'b01111; w[119][119] = 5'b00000; w[119][120] = 5'b10000; w[119][121] = 5'b10000; w[119][122] = 5'b10000; w[119][123] = 5'b10000; w[119][124] = 5'b10000; w[119][125] = 5'b10000; w[119][126] = 5'b10000; w[119][127] = 5'b10000; w[119][128] = 5'b10000; w[119][129] = 5'b10000; w[119][130] = 5'b00000; w[119][131] = 5'b10000; w[119][132] = 5'b01111; w[119][133] = 5'b01111; w[119][134] = 5'b00000; w[119][135] = 5'b00000; w[119][136] = 5'b10000; w[119][137] = 5'b10000; w[119][138] = 5'b10000; w[119][139] = 5'b10000; w[119][140] = 5'b10000; w[119][141] = 5'b10000; w[119][142] = 5'b10000; w[119][143] = 5'b10000; w[119][144] = 5'b10000; w[119][145] = 5'b10000; w[119][146] = 5'b01111; w[119][147] = 5'b01111; w[119][148] = 5'b00000; w[119][149] = 5'b10000; w[119][150] = 5'b10000; w[119][151] = 5'b10000; w[119][152] = 5'b10000; w[119][153] = 5'b10000; w[119][154] = 5'b10000; w[119][155] = 5'b10000; w[119][156] = 5'b10000; w[119][157] = 5'b10000; w[119][158] = 5'b10000; w[119][159] = 5'b10000; w[119][160] = 5'b00000; w[119][161] = 5'b00000; w[119][162] = 5'b00000; w[119][163] = 5'b10000; w[119][164] = 5'b10000; w[119][165] = 5'b10000; w[119][166] = 5'b10000; w[119][167] = 5'b10000; w[119][168] = 5'b10000; w[119][169] = 5'b10000; w[119][170] = 5'b10000; w[119][171] = 5'b00000; w[119][172] = 5'b10000; w[119][173] = 5'b10000; w[119][174] = 5'b00000; w[119][175] = 5'b00000; w[119][176] = 5'b00000; w[119][177] = 5'b10000; w[119][178] = 5'b00000; w[119][179] = 5'b10000; w[119][180] = 5'b10000; w[119][181] = 5'b10000; w[119][182] = 5'b10000; w[119][183] = 5'b10000; w[119][184] = 5'b10000; w[119][185] = 5'b10000; w[119][186] = 5'b10000; w[119][187] = 5'b10000; w[119][188] = 5'b10000; w[119][189] = 5'b10000; w[119][190] = 5'b10000; w[119][191] = 5'b10000; w[119][192] = 5'b10000; w[119][193] = 5'b10000; w[119][194] = 5'b10000; w[119][195] = 5'b10000; w[119][196] = 5'b10000; w[119][197] = 5'b10000; w[119][198] = 5'b10000; w[119][199] = 5'b10000; w[119][200] = 5'b10000; w[119][201] = 5'b10000; w[119][202] = 5'b10000; w[119][203] = 5'b10000; w[119][204] = 5'b10000; w[119][205] = 5'b10000; w[119][206] = 5'b10000; w[119][207] = 5'b10000; w[119][208] = 5'b10000; w[119][209] = 5'b10000; 
w[120][0] = 5'b00000; w[120][1] = 5'b00000; w[120][2] = 5'b00000; w[120][3] = 5'b00000; w[120][4] = 5'b00000; w[120][5] = 5'b00000; w[120][6] = 5'b00000; w[120][7] = 5'b00000; w[120][8] = 5'b00000; w[120][9] = 5'b00000; w[120][10] = 5'b00000; w[120][11] = 5'b00000; w[120][12] = 5'b00000; w[120][13] = 5'b00000; w[120][14] = 5'b00000; w[120][15] = 5'b00000; w[120][16] = 5'b00000; w[120][17] = 5'b00000; w[120][18] = 5'b00000; w[120][19] = 5'b00000; w[120][20] = 5'b00000; w[120][21] = 5'b00000; w[120][22] = 5'b00000; w[120][23] = 5'b00000; w[120][24] = 5'b00000; w[120][25] = 5'b00000; w[120][26] = 5'b00000; w[120][27] = 5'b00000; w[120][28] = 5'b00000; w[120][29] = 5'b00000; w[120][30] = 5'b10000; w[120][31] = 5'b00000; w[120][32] = 5'b01111; w[120][33] = 5'b00000; w[120][34] = 5'b10000; w[120][35] = 5'b10000; w[120][36] = 5'b10000; w[120][37] = 5'b01111; w[120][38] = 5'b00000; w[120][39] = 5'b10000; w[120][40] = 5'b00000; w[120][41] = 5'b00000; w[120][42] = 5'b00000; w[120][43] = 5'b00000; w[120][44] = 5'b10000; w[120][45] = 5'b01111; w[120][46] = 5'b01111; w[120][47] = 5'b00000; w[120][48] = 5'b10000; w[120][49] = 5'b10000; w[120][50] = 5'b10000; w[120][51] = 5'b01111; w[120][52] = 5'b01111; w[120][53] = 5'b10000; w[120][54] = 5'b00000; w[120][55] = 5'b00000; w[120][56] = 5'b00000; w[120][57] = 5'b00000; w[120][58] = 5'b01111; w[120][59] = 5'b01111; w[120][60] = 5'b01111; w[120][61] = 5'b01111; w[120][62] = 5'b10000; w[120][63] = 5'b10000; w[120][64] = 5'b00000; w[120][65] = 5'b01111; w[120][66] = 5'b01111; w[120][67] = 5'b01111; w[120][68] = 5'b00000; w[120][69] = 5'b00000; w[120][70] = 5'b00000; w[120][71] = 5'b00000; w[120][72] = 5'b01111; w[120][73] = 5'b01111; w[120][74] = 5'b01111; w[120][75] = 5'b01111; w[120][76] = 5'b10000; w[120][77] = 5'b10000; w[120][78] = 5'b00000; w[120][79] = 5'b01111; w[120][80] = 5'b01111; w[120][81] = 5'b01111; w[120][82] = 5'b00000; w[120][83] = 5'b00000; w[120][84] = 5'b00000; w[120][85] = 5'b00000; w[120][86] = 5'b01111; w[120][87] = 5'b01111; w[120][88] = 5'b01111; w[120][89] = 5'b01111; w[120][90] = 5'b10000; w[120][91] = 5'b10000; w[120][92] = 5'b00000; w[120][93] = 5'b01111; w[120][94] = 5'b01111; w[120][95] = 5'b00000; w[120][96] = 5'b00000; w[120][97] = 5'b00000; w[120][98] = 5'b00000; w[120][99] = 5'b00000; w[120][100] = 5'b01111; w[120][101] = 5'b01111; w[120][102] = 5'b01111; w[120][103] = 5'b00000; w[120][104] = 5'b10000; w[120][105] = 5'b10000; w[120][106] = 5'b01111; w[120][107] = 5'b01111; w[120][108] = 5'b01111; w[120][109] = 5'b01111; w[120][110] = 5'b00000; w[120][111] = 5'b00000; w[120][112] = 5'b00000; w[120][113] = 5'b00000; w[120][114] = 5'b01111; w[120][115] = 5'b01111; w[120][116] = 5'b01111; w[120][117] = 5'b00000; w[120][118] = 5'b10000; w[120][119] = 5'b10000; w[120][120] = 5'b00000; w[120][121] = 5'b01111; w[120][122] = 5'b01111; w[120][123] = 5'b01111; w[120][124] = 5'b00000; w[120][125] = 5'b00000; w[120][126] = 5'b00000; w[120][127] = 5'b00000; w[120][128] = 5'b01111; w[120][129] = 5'b01111; w[120][130] = 5'b01111; w[120][131] = 5'b00000; w[120][132] = 5'b10000; w[120][133] = 5'b10000; w[120][134] = 5'b01111; w[120][135] = 5'b01111; w[120][136] = 5'b01111; w[120][137] = 5'b01111; w[120][138] = 5'b00000; w[120][139] = 5'b00000; w[120][140] = 5'b00000; w[120][141] = 5'b00000; w[120][142] = 5'b01111; w[120][143] = 5'b01111; w[120][144] = 5'b01111; w[120][145] = 5'b00000; w[120][146] = 5'b10000; w[120][147] = 5'b10000; w[120][148] = 5'b01111; w[120][149] = 5'b01111; w[120][150] = 5'b01111; w[120][151] = 5'b01111; w[120][152] = 5'b00000; w[120][153] = 5'b00000; w[120][154] = 5'b00000; w[120][155] = 5'b00000; w[120][156] = 5'b00000; w[120][157] = 5'b01111; w[120][158] = 5'b01111; w[120][159] = 5'b00000; w[120][160] = 5'b10000; w[120][161] = 5'b10000; w[120][162] = 5'b01111; w[120][163] = 5'b01111; w[120][164] = 5'b01111; w[120][165] = 5'b00000; w[120][166] = 5'b00000; w[120][167] = 5'b00000; w[120][168] = 5'b00000; w[120][169] = 5'b00000; w[120][170] = 5'b00000; w[120][171] = 5'b01111; w[120][172] = 5'b01111; w[120][173] = 5'b00000; w[120][174] = 5'b10000; w[120][175] = 5'b10000; w[120][176] = 5'b01111; w[120][177] = 5'b01111; w[120][178] = 5'b01111; w[120][179] = 5'b00000; w[120][180] = 5'b00000; w[120][181] = 5'b00000; w[120][182] = 5'b00000; w[120][183] = 5'b00000; w[120][184] = 5'b00000; w[120][185] = 5'b00000; w[120][186] = 5'b00000; w[120][187] = 5'b00000; w[120][188] = 5'b00000; w[120][189] = 5'b00000; w[120][190] = 5'b00000; w[120][191] = 5'b00000; w[120][192] = 5'b00000; w[120][193] = 5'b00000; w[120][194] = 5'b00000; w[120][195] = 5'b00000; w[120][196] = 5'b00000; w[120][197] = 5'b00000; w[120][198] = 5'b00000; w[120][199] = 5'b00000; w[120][200] = 5'b00000; w[120][201] = 5'b00000; w[120][202] = 5'b00000; w[120][203] = 5'b00000; w[120][204] = 5'b00000; w[120][205] = 5'b00000; w[120][206] = 5'b00000; w[120][207] = 5'b00000; w[120][208] = 5'b00000; w[120][209] = 5'b00000; 
w[121][0] = 5'b00000; w[121][1] = 5'b00000; w[121][2] = 5'b00000; w[121][3] = 5'b00000; w[121][4] = 5'b00000; w[121][5] = 5'b00000; w[121][6] = 5'b00000; w[121][7] = 5'b00000; w[121][8] = 5'b00000; w[121][9] = 5'b00000; w[121][10] = 5'b00000; w[121][11] = 5'b00000; w[121][12] = 5'b00000; w[121][13] = 5'b00000; w[121][14] = 5'b00000; w[121][15] = 5'b00000; w[121][16] = 5'b00000; w[121][17] = 5'b00000; w[121][18] = 5'b00000; w[121][19] = 5'b00000; w[121][20] = 5'b00000; w[121][21] = 5'b00000; w[121][22] = 5'b00000; w[121][23] = 5'b00000; w[121][24] = 5'b00000; w[121][25] = 5'b00000; w[121][26] = 5'b00000; w[121][27] = 5'b00000; w[121][28] = 5'b00000; w[121][29] = 5'b00000; w[121][30] = 5'b10000; w[121][31] = 5'b00000; w[121][32] = 5'b01111; w[121][33] = 5'b00000; w[121][34] = 5'b10000; w[121][35] = 5'b10000; w[121][36] = 5'b10000; w[121][37] = 5'b01111; w[121][38] = 5'b00000; w[121][39] = 5'b10000; w[121][40] = 5'b00000; w[121][41] = 5'b00000; w[121][42] = 5'b00000; w[121][43] = 5'b00000; w[121][44] = 5'b10000; w[121][45] = 5'b01111; w[121][46] = 5'b01111; w[121][47] = 5'b00000; w[121][48] = 5'b10000; w[121][49] = 5'b10000; w[121][50] = 5'b10000; w[121][51] = 5'b01111; w[121][52] = 5'b01111; w[121][53] = 5'b10000; w[121][54] = 5'b00000; w[121][55] = 5'b00000; w[121][56] = 5'b00000; w[121][57] = 5'b00000; w[121][58] = 5'b01111; w[121][59] = 5'b01111; w[121][60] = 5'b01111; w[121][61] = 5'b01111; w[121][62] = 5'b10000; w[121][63] = 5'b10000; w[121][64] = 5'b00000; w[121][65] = 5'b01111; w[121][66] = 5'b01111; w[121][67] = 5'b01111; w[121][68] = 5'b00000; w[121][69] = 5'b00000; w[121][70] = 5'b00000; w[121][71] = 5'b00000; w[121][72] = 5'b01111; w[121][73] = 5'b01111; w[121][74] = 5'b01111; w[121][75] = 5'b01111; w[121][76] = 5'b10000; w[121][77] = 5'b10000; w[121][78] = 5'b00000; w[121][79] = 5'b01111; w[121][80] = 5'b01111; w[121][81] = 5'b01111; w[121][82] = 5'b00000; w[121][83] = 5'b00000; w[121][84] = 5'b00000; w[121][85] = 5'b00000; w[121][86] = 5'b01111; w[121][87] = 5'b01111; w[121][88] = 5'b01111; w[121][89] = 5'b01111; w[121][90] = 5'b10000; w[121][91] = 5'b10000; w[121][92] = 5'b00000; w[121][93] = 5'b01111; w[121][94] = 5'b01111; w[121][95] = 5'b00000; w[121][96] = 5'b00000; w[121][97] = 5'b00000; w[121][98] = 5'b00000; w[121][99] = 5'b00000; w[121][100] = 5'b01111; w[121][101] = 5'b01111; w[121][102] = 5'b01111; w[121][103] = 5'b00000; w[121][104] = 5'b10000; w[121][105] = 5'b10000; w[121][106] = 5'b01111; w[121][107] = 5'b01111; w[121][108] = 5'b01111; w[121][109] = 5'b01111; w[121][110] = 5'b00000; w[121][111] = 5'b00000; w[121][112] = 5'b00000; w[121][113] = 5'b00000; w[121][114] = 5'b01111; w[121][115] = 5'b01111; w[121][116] = 5'b01111; w[121][117] = 5'b00000; w[121][118] = 5'b10000; w[121][119] = 5'b10000; w[121][120] = 5'b01111; w[121][121] = 5'b00000; w[121][122] = 5'b01111; w[121][123] = 5'b01111; w[121][124] = 5'b00000; w[121][125] = 5'b00000; w[121][126] = 5'b00000; w[121][127] = 5'b00000; w[121][128] = 5'b01111; w[121][129] = 5'b01111; w[121][130] = 5'b01111; w[121][131] = 5'b00000; w[121][132] = 5'b10000; w[121][133] = 5'b10000; w[121][134] = 5'b01111; w[121][135] = 5'b01111; w[121][136] = 5'b01111; w[121][137] = 5'b01111; w[121][138] = 5'b00000; w[121][139] = 5'b00000; w[121][140] = 5'b00000; w[121][141] = 5'b00000; w[121][142] = 5'b01111; w[121][143] = 5'b01111; w[121][144] = 5'b01111; w[121][145] = 5'b00000; w[121][146] = 5'b10000; w[121][147] = 5'b10000; w[121][148] = 5'b01111; w[121][149] = 5'b01111; w[121][150] = 5'b01111; w[121][151] = 5'b01111; w[121][152] = 5'b00000; w[121][153] = 5'b00000; w[121][154] = 5'b00000; w[121][155] = 5'b00000; w[121][156] = 5'b00000; w[121][157] = 5'b01111; w[121][158] = 5'b01111; w[121][159] = 5'b00000; w[121][160] = 5'b10000; w[121][161] = 5'b10000; w[121][162] = 5'b01111; w[121][163] = 5'b01111; w[121][164] = 5'b01111; w[121][165] = 5'b00000; w[121][166] = 5'b00000; w[121][167] = 5'b00000; w[121][168] = 5'b00000; w[121][169] = 5'b00000; w[121][170] = 5'b00000; w[121][171] = 5'b01111; w[121][172] = 5'b01111; w[121][173] = 5'b00000; w[121][174] = 5'b10000; w[121][175] = 5'b10000; w[121][176] = 5'b01111; w[121][177] = 5'b01111; w[121][178] = 5'b01111; w[121][179] = 5'b00000; w[121][180] = 5'b00000; w[121][181] = 5'b00000; w[121][182] = 5'b00000; w[121][183] = 5'b00000; w[121][184] = 5'b00000; w[121][185] = 5'b00000; w[121][186] = 5'b00000; w[121][187] = 5'b00000; w[121][188] = 5'b00000; w[121][189] = 5'b00000; w[121][190] = 5'b00000; w[121][191] = 5'b00000; w[121][192] = 5'b00000; w[121][193] = 5'b00000; w[121][194] = 5'b00000; w[121][195] = 5'b00000; w[121][196] = 5'b00000; w[121][197] = 5'b00000; w[121][198] = 5'b00000; w[121][199] = 5'b00000; w[121][200] = 5'b00000; w[121][201] = 5'b00000; w[121][202] = 5'b00000; w[121][203] = 5'b00000; w[121][204] = 5'b00000; w[121][205] = 5'b00000; w[121][206] = 5'b00000; w[121][207] = 5'b00000; w[121][208] = 5'b00000; w[121][209] = 5'b00000; 
w[122][0] = 5'b00000; w[122][1] = 5'b00000; w[122][2] = 5'b00000; w[122][3] = 5'b00000; w[122][4] = 5'b00000; w[122][5] = 5'b00000; w[122][6] = 5'b00000; w[122][7] = 5'b00000; w[122][8] = 5'b00000; w[122][9] = 5'b00000; w[122][10] = 5'b00000; w[122][11] = 5'b00000; w[122][12] = 5'b00000; w[122][13] = 5'b00000; w[122][14] = 5'b00000; w[122][15] = 5'b00000; w[122][16] = 5'b00000; w[122][17] = 5'b00000; w[122][18] = 5'b00000; w[122][19] = 5'b00000; w[122][20] = 5'b00000; w[122][21] = 5'b00000; w[122][22] = 5'b00000; w[122][23] = 5'b00000; w[122][24] = 5'b00000; w[122][25] = 5'b00000; w[122][26] = 5'b00000; w[122][27] = 5'b00000; w[122][28] = 5'b00000; w[122][29] = 5'b00000; w[122][30] = 5'b10000; w[122][31] = 5'b00000; w[122][32] = 5'b01111; w[122][33] = 5'b00000; w[122][34] = 5'b10000; w[122][35] = 5'b10000; w[122][36] = 5'b10000; w[122][37] = 5'b01111; w[122][38] = 5'b00000; w[122][39] = 5'b10000; w[122][40] = 5'b00000; w[122][41] = 5'b00000; w[122][42] = 5'b00000; w[122][43] = 5'b00000; w[122][44] = 5'b10000; w[122][45] = 5'b01111; w[122][46] = 5'b01111; w[122][47] = 5'b00000; w[122][48] = 5'b10000; w[122][49] = 5'b10000; w[122][50] = 5'b10000; w[122][51] = 5'b01111; w[122][52] = 5'b01111; w[122][53] = 5'b10000; w[122][54] = 5'b00000; w[122][55] = 5'b00000; w[122][56] = 5'b00000; w[122][57] = 5'b00000; w[122][58] = 5'b01111; w[122][59] = 5'b01111; w[122][60] = 5'b01111; w[122][61] = 5'b01111; w[122][62] = 5'b10000; w[122][63] = 5'b10000; w[122][64] = 5'b00000; w[122][65] = 5'b01111; w[122][66] = 5'b01111; w[122][67] = 5'b01111; w[122][68] = 5'b00000; w[122][69] = 5'b00000; w[122][70] = 5'b00000; w[122][71] = 5'b00000; w[122][72] = 5'b01111; w[122][73] = 5'b01111; w[122][74] = 5'b01111; w[122][75] = 5'b01111; w[122][76] = 5'b10000; w[122][77] = 5'b10000; w[122][78] = 5'b00000; w[122][79] = 5'b01111; w[122][80] = 5'b01111; w[122][81] = 5'b01111; w[122][82] = 5'b00000; w[122][83] = 5'b00000; w[122][84] = 5'b00000; w[122][85] = 5'b00000; w[122][86] = 5'b01111; w[122][87] = 5'b01111; w[122][88] = 5'b01111; w[122][89] = 5'b01111; w[122][90] = 5'b10000; w[122][91] = 5'b10000; w[122][92] = 5'b00000; w[122][93] = 5'b01111; w[122][94] = 5'b01111; w[122][95] = 5'b00000; w[122][96] = 5'b00000; w[122][97] = 5'b00000; w[122][98] = 5'b00000; w[122][99] = 5'b00000; w[122][100] = 5'b01111; w[122][101] = 5'b01111; w[122][102] = 5'b01111; w[122][103] = 5'b00000; w[122][104] = 5'b10000; w[122][105] = 5'b10000; w[122][106] = 5'b01111; w[122][107] = 5'b01111; w[122][108] = 5'b01111; w[122][109] = 5'b01111; w[122][110] = 5'b00000; w[122][111] = 5'b00000; w[122][112] = 5'b00000; w[122][113] = 5'b00000; w[122][114] = 5'b01111; w[122][115] = 5'b01111; w[122][116] = 5'b01111; w[122][117] = 5'b00000; w[122][118] = 5'b10000; w[122][119] = 5'b10000; w[122][120] = 5'b01111; w[122][121] = 5'b01111; w[122][122] = 5'b00000; w[122][123] = 5'b01111; w[122][124] = 5'b00000; w[122][125] = 5'b00000; w[122][126] = 5'b00000; w[122][127] = 5'b00000; w[122][128] = 5'b01111; w[122][129] = 5'b01111; w[122][130] = 5'b01111; w[122][131] = 5'b00000; w[122][132] = 5'b10000; w[122][133] = 5'b10000; w[122][134] = 5'b01111; w[122][135] = 5'b01111; w[122][136] = 5'b01111; w[122][137] = 5'b01111; w[122][138] = 5'b00000; w[122][139] = 5'b00000; w[122][140] = 5'b00000; w[122][141] = 5'b00000; w[122][142] = 5'b01111; w[122][143] = 5'b01111; w[122][144] = 5'b01111; w[122][145] = 5'b00000; w[122][146] = 5'b10000; w[122][147] = 5'b10000; w[122][148] = 5'b01111; w[122][149] = 5'b01111; w[122][150] = 5'b01111; w[122][151] = 5'b01111; w[122][152] = 5'b00000; w[122][153] = 5'b00000; w[122][154] = 5'b00000; w[122][155] = 5'b00000; w[122][156] = 5'b00000; w[122][157] = 5'b01111; w[122][158] = 5'b01111; w[122][159] = 5'b00000; w[122][160] = 5'b10000; w[122][161] = 5'b10000; w[122][162] = 5'b01111; w[122][163] = 5'b01111; w[122][164] = 5'b01111; w[122][165] = 5'b00000; w[122][166] = 5'b00000; w[122][167] = 5'b00000; w[122][168] = 5'b00000; w[122][169] = 5'b00000; w[122][170] = 5'b00000; w[122][171] = 5'b01111; w[122][172] = 5'b01111; w[122][173] = 5'b00000; w[122][174] = 5'b10000; w[122][175] = 5'b10000; w[122][176] = 5'b01111; w[122][177] = 5'b01111; w[122][178] = 5'b01111; w[122][179] = 5'b00000; w[122][180] = 5'b00000; w[122][181] = 5'b00000; w[122][182] = 5'b00000; w[122][183] = 5'b00000; w[122][184] = 5'b00000; w[122][185] = 5'b00000; w[122][186] = 5'b00000; w[122][187] = 5'b00000; w[122][188] = 5'b00000; w[122][189] = 5'b00000; w[122][190] = 5'b00000; w[122][191] = 5'b00000; w[122][192] = 5'b00000; w[122][193] = 5'b00000; w[122][194] = 5'b00000; w[122][195] = 5'b00000; w[122][196] = 5'b00000; w[122][197] = 5'b00000; w[122][198] = 5'b00000; w[122][199] = 5'b00000; w[122][200] = 5'b00000; w[122][201] = 5'b00000; w[122][202] = 5'b00000; w[122][203] = 5'b00000; w[122][204] = 5'b00000; w[122][205] = 5'b00000; w[122][206] = 5'b00000; w[122][207] = 5'b00000; w[122][208] = 5'b00000; w[122][209] = 5'b00000; 
w[123][0] = 5'b01111; w[123][1] = 5'b01111; w[123][2] = 5'b01111; w[123][3] = 5'b01111; w[123][4] = 5'b01111; w[123][5] = 5'b01111; w[123][6] = 5'b01111; w[123][7] = 5'b01111; w[123][8] = 5'b01111; w[123][9] = 5'b01111; w[123][10] = 5'b01111; w[123][11] = 5'b01111; w[123][12] = 5'b01111; w[123][13] = 5'b01111; w[123][14] = 5'b01111; w[123][15] = 5'b01111; w[123][16] = 5'b01111; w[123][17] = 5'b01111; w[123][18] = 5'b01111; w[123][19] = 5'b01111; w[123][20] = 5'b01111; w[123][21] = 5'b01111; w[123][22] = 5'b01111; w[123][23] = 5'b01111; w[123][24] = 5'b01111; w[123][25] = 5'b01111; w[123][26] = 5'b01111; w[123][27] = 5'b01111; w[123][28] = 5'b01111; w[123][29] = 5'b01111; w[123][30] = 5'b00000; w[123][31] = 5'b10000; w[123][32] = 5'b00000; w[123][33] = 5'b10000; w[123][34] = 5'b00000; w[123][35] = 5'b00000; w[123][36] = 5'b00000; w[123][37] = 5'b00000; w[123][38] = 5'b10000; w[123][39] = 5'b00000; w[123][40] = 5'b01111; w[123][41] = 5'b01111; w[123][42] = 5'b01111; w[123][43] = 5'b01111; w[123][44] = 5'b00000; w[123][45] = 5'b00000; w[123][46] = 5'b00000; w[123][47] = 5'b10000; w[123][48] = 5'b00000; w[123][49] = 5'b00000; w[123][50] = 5'b00000; w[123][51] = 5'b00000; w[123][52] = 5'b00000; w[123][53] = 5'b00000; w[123][54] = 5'b01111; w[123][55] = 5'b01111; w[123][56] = 5'b01111; w[123][57] = 5'b01111; w[123][58] = 5'b01111; w[123][59] = 5'b01111; w[123][60] = 5'b01111; w[123][61] = 5'b00000; w[123][62] = 5'b10000; w[123][63] = 5'b10000; w[123][64] = 5'b01111; w[123][65] = 5'b01111; w[123][66] = 5'b01111; w[123][67] = 5'b01111; w[123][68] = 5'b01111; w[123][69] = 5'b01111; w[123][70] = 5'b01111; w[123][71] = 5'b01111; w[123][72] = 5'b01111; w[123][73] = 5'b01111; w[123][74] = 5'b00000; w[123][75] = 5'b00000; w[123][76] = 5'b10000; w[123][77] = 5'b10000; w[123][78] = 5'b01111; w[123][79] = 5'b00000; w[123][80] = 5'b01111; w[123][81] = 5'b01111; w[123][82] = 5'b01111; w[123][83] = 5'b01111; w[123][84] = 5'b01111; w[123][85] = 5'b01111; w[123][86] = 5'b01111; w[123][87] = 5'b01111; w[123][88] = 5'b00000; w[123][89] = 5'b00000; w[123][90] = 5'b10000; w[123][91] = 5'b10000; w[123][92] = 5'b01111; w[123][93] = 5'b00000; w[123][94] = 5'b00000; w[123][95] = 5'b01111; w[123][96] = 5'b01111; w[123][97] = 5'b01111; w[123][98] = 5'b01111; w[123][99] = 5'b01111; w[123][100] = 5'b01111; w[123][101] = 5'b01111; w[123][102] = 5'b00000; w[123][103] = 5'b01111; w[123][104] = 5'b10000; w[123][105] = 5'b10000; w[123][106] = 5'b01111; w[123][107] = 5'b01111; w[123][108] = 5'b01111; w[123][109] = 5'b01111; w[123][110] = 5'b01111; w[123][111] = 5'b01111; w[123][112] = 5'b01111; w[123][113] = 5'b01111; w[123][114] = 5'b01111; w[123][115] = 5'b01111; w[123][116] = 5'b00000; w[123][117] = 5'b01111; w[123][118] = 5'b10000; w[123][119] = 5'b10000; w[123][120] = 5'b01111; w[123][121] = 5'b01111; w[123][122] = 5'b01111; w[123][123] = 5'b00000; w[123][124] = 5'b01111; w[123][125] = 5'b01111; w[123][126] = 5'b01111; w[123][127] = 5'b01111; w[123][128] = 5'b01111; w[123][129] = 5'b01111; w[123][130] = 5'b00000; w[123][131] = 5'b01111; w[123][132] = 5'b10000; w[123][133] = 5'b10000; w[123][134] = 5'b00000; w[123][135] = 5'b00000; w[123][136] = 5'b01111; w[123][137] = 5'b01111; w[123][138] = 5'b01111; w[123][139] = 5'b01111; w[123][140] = 5'b01111; w[123][141] = 5'b01111; w[123][142] = 5'b01111; w[123][143] = 5'b01111; w[123][144] = 5'b01111; w[123][145] = 5'b01111; w[123][146] = 5'b10000; w[123][147] = 5'b10000; w[123][148] = 5'b00000; w[123][149] = 5'b01111; w[123][150] = 5'b01111; w[123][151] = 5'b01111; w[123][152] = 5'b01111; w[123][153] = 5'b01111; w[123][154] = 5'b01111; w[123][155] = 5'b01111; w[123][156] = 5'b01111; w[123][157] = 5'b01111; w[123][158] = 5'b01111; w[123][159] = 5'b01111; w[123][160] = 5'b00000; w[123][161] = 5'b00000; w[123][162] = 5'b00000; w[123][163] = 5'b01111; w[123][164] = 5'b01111; w[123][165] = 5'b01111; w[123][166] = 5'b01111; w[123][167] = 5'b01111; w[123][168] = 5'b01111; w[123][169] = 5'b01111; w[123][170] = 5'b01111; w[123][171] = 5'b00000; w[123][172] = 5'b01111; w[123][173] = 5'b01111; w[123][174] = 5'b00000; w[123][175] = 5'b00000; w[123][176] = 5'b00000; w[123][177] = 5'b01111; w[123][178] = 5'b00000; w[123][179] = 5'b01111; w[123][180] = 5'b01111; w[123][181] = 5'b01111; w[123][182] = 5'b01111; w[123][183] = 5'b01111; w[123][184] = 5'b01111; w[123][185] = 5'b01111; w[123][186] = 5'b01111; w[123][187] = 5'b01111; w[123][188] = 5'b01111; w[123][189] = 5'b01111; w[123][190] = 5'b01111; w[123][191] = 5'b01111; w[123][192] = 5'b01111; w[123][193] = 5'b01111; w[123][194] = 5'b01111; w[123][195] = 5'b01111; w[123][196] = 5'b01111; w[123][197] = 5'b01111; w[123][198] = 5'b01111; w[123][199] = 5'b01111; w[123][200] = 5'b01111; w[123][201] = 5'b01111; w[123][202] = 5'b01111; w[123][203] = 5'b01111; w[123][204] = 5'b01111; w[123][205] = 5'b01111; w[123][206] = 5'b01111; w[123][207] = 5'b01111; w[123][208] = 5'b01111; w[123][209] = 5'b01111; 
w[124][0] = 5'b01111; w[124][1] = 5'b01111; w[124][2] = 5'b01111; w[124][3] = 5'b01111; w[124][4] = 5'b01111; w[124][5] = 5'b01111; w[124][6] = 5'b01111; w[124][7] = 5'b01111; w[124][8] = 5'b01111; w[124][9] = 5'b01111; w[124][10] = 5'b01111; w[124][11] = 5'b01111; w[124][12] = 5'b01111; w[124][13] = 5'b01111; w[124][14] = 5'b01111; w[124][15] = 5'b01111; w[124][16] = 5'b01111; w[124][17] = 5'b01111; w[124][18] = 5'b01111; w[124][19] = 5'b01111; w[124][20] = 5'b01111; w[124][21] = 5'b01111; w[124][22] = 5'b01111; w[124][23] = 5'b01111; w[124][24] = 5'b01111; w[124][25] = 5'b01111; w[124][26] = 5'b01111; w[124][27] = 5'b01111; w[124][28] = 5'b01111; w[124][29] = 5'b01111; w[124][30] = 5'b01111; w[124][31] = 5'b00000; w[124][32] = 5'b10000; w[124][33] = 5'b10000; w[124][34] = 5'b10000; w[124][35] = 5'b10000; w[124][36] = 5'b10000; w[124][37] = 5'b10000; w[124][38] = 5'b00000; w[124][39] = 5'b01111; w[124][40] = 5'b01111; w[124][41] = 5'b01111; w[124][42] = 5'b01111; w[124][43] = 5'b01111; w[124][44] = 5'b01111; w[124][45] = 5'b10000; w[124][46] = 5'b10000; w[124][47] = 5'b10000; w[124][48] = 5'b10000; w[124][49] = 5'b10000; w[124][50] = 5'b10000; w[124][51] = 5'b10000; w[124][52] = 5'b10000; w[124][53] = 5'b01111; w[124][54] = 5'b01111; w[124][55] = 5'b01111; w[124][56] = 5'b01111; w[124][57] = 5'b01111; w[124][58] = 5'b01111; w[124][59] = 5'b00000; w[124][60] = 5'b00000; w[124][61] = 5'b01111; w[124][62] = 5'b10000; w[124][63] = 5'b00000; w[124][64] = 5'b01111; w[124][65] = 5'b00000; w[124][66] = 5'b00000; w[124][67] = 5'b01111; w[124][68] = 5'b01111; w[124][69] = 5'b01111; w[124][70] = 5'b01111; w[124][71] = 5'b01111; w[124][72] = 5'b01111; w[124][73] = 5'b00000; w[124][74] = 5'b01111; w[124][75] = 5'b01111; w[124][76] = 5'b10000; w[124][77] = 5'b00000; w[124][78] = 5'b01111; w[124][79] = 5'b01111; w[124][80] = 5'b00000; w[124][81] = 5'b01111; w[124][82] = 5'b01111; w[124][83] = 5'b01111; w[124][84] = 5'b01111; w[124][85] = 5'b01111; w[124][86] = 5'b01111; w[124][87] = 5'b00000; w[124][88] = 5'b01111; w[124][89] = 5'b01111; w[124][90] = 5'b10000; w[124][91] = 5'b10000; w[124][92] = 5'b01111; w[124][93] = 5'b01111; w[124][94] = 5'b01111; w[124][95] = 5'b01111; w[124][96] = 5'b01111; w[124][97] = 5'b01111; w[124][98] = 5'b01111; w[124][99] = 5'b01111; w[124][100] = 5'b01111; w[124][101] = 5'b00000; w[124][102] = 5'b01111; w[124][103] = 5'b01111; w[124][104] = 5'b10000; w[124][105] = 5'b10000; w[124][106] = 5'b01111; w[124][107] = 5'b00000; w[124][108] = 5'b00000; w[124][109] = 5'b01111; w[124][110] = 5'b01111; w[124][111] = 5'b01111; w[124][112] = 5'b01111; w[124][113] = 5'b01111; w[124][114] = 5'b01111; w[124][115] = 5'b00000; w[124][116] = 5'b01111; w[124][117] = 5'b01111; w[124][118] = 5'b10000; w[124][119] = 5'b10000; w[124][120] = 5'b00000; w[124][121] = 5'b00000; w[124][122] = 5'b00000; w[124][123] = 5'b01111; w[124][124] = 5'b00000; w[124][125] = 5'b01111; w[124][126] = 5'b01111; w[124][127] = 5'b01111; w[124][128] = 5'b01111; w[124][129] = 5'b00000; w[124][130] = 5'b01111; w[124][131] = 5'b01111; w[124][132] = 5'b00000; w[124][133] = 5'b10000; w[124][134] = 5'b01111; w[124][135] = 5'b01111; w[124][136] = 5'b00000; w[124][137] = 5'b01111; w[124][138] = 5'b01111; w[124][139] = 5'b01111; w[124][140] = 5'b01111; w[124][141] = 5'b01111; w[124][142] = 5'b01111; w[124][143] = 5'b00000; w[124][144] = 5'b00000; w[124][145] = 5'b01111; w[124][146] = 5'b00000; w[124][147] = 5'b10000; w[124][148] = 5'b01111; w[124][149] = 5'b00000; w[124][150] = 5'b00000; w[124][151] = 5'b01111; w[124][152] = 5'b01111; w[124][153] = 5'b01111; w[124][154] = 5'b01111; w[124][155] = 5'b01111; w[124][156] = 5'b01111; w[124][157] = 5'b00000; w[124][158] = 5'b00000; w[124][159] = 5'b00000; w[124][160] = 5'b10000; w[124][161] = 5'b10000; w[124][162] = 5'b10000; w[124][163] = 5'b00000; w[124][164] = 5'b00000; w[124][165] = 5'b01111; w[124][166] = 5'b01111; w[124][167] = 5'b01111; w[124][168] = 5'b01111; w[124][169] = 5'b01111; w[124][170] = 5'b01111; w[124][171] = 5'b01111; w[124][172] = 5'b00000; w[124][173] = 5'b00000; w[124][174] = 5'b10000; w[124][175] = 5'b10000; w[124][176] = 5'b10000; w[124][177] = 5'b00000; w[124][178] = 5'b01111; w[124][179] = 5'b01111; w[124][180] = 5'b01111; w[124][181] = 5'b01111; w[124][182] = 5'b01111; w[124][183] = 5'b01111; w[124][184] = 5'b01111; w[124][185] = 5'b01111; w[124][186] = 5'b01111; w[124][187] = 5'b01111; w[124][188] = 5'b01111; w[124][189] = 5'b01111; w[124][190] = 5'b01111; w[124][191] = 5'b01111; w[124][192] = 5'b01111; w[124][193] = 5'b01111; w[124][194] = 5'b01111; w[124][195] = 5'b01111; w[124][196] = 5'b01111; w[124][197] = 5'b01111; w[124][198] = 5'b01111; w[124][199] = 5'b01111; w[124][200] = 5'b01111; w[124][201] = 5'b01111; w[124][202] = 5'b01111; w[124][203] = 5'b01111; w[124][204] = 5'b01111; w[124][205] = 5'b01111; w[124][206] = 5'b01111; w[124][207] = 5'b01111; w[124][208] = 5'b01111; w[124][209] = 5'b01111; 
w[125][0] = 5'b01111; w[125][1] = 5'b01111; w[125][2] = 5'b01111; w[125][3] = 5'b01111; w[125][4] = 5'b01111; w[125][5] = 5'b01111; w[125][6] = 5'b01111; w[125][7] = 5'b01111; w[125][8] = 5'b01111; w[125][9] = 5'b01111; w[125][10] = 5'b01111; w[125][11] = 5'b01111; w[125][12] = 5'b01111; w[125][13] = 5'b01111; w[125][14] = 5'b01111; w[125][15] = 5'b01111; w[125][16] = 5'b01111; w[125][17] = 5'b01111; w[125][18] = 5'b01111; w[125][19] = 5'b01111; w[125][20] = 5'b01111; w[125][21] = 5'b01111; w[125][22] = 5'b01111; w[125][23] = 5'b01111; w[125][24] = 5'b01111; w[125][25] = 5'b01111; w[125][26] = 5'b01111; w[125][27] = 5'b01111; w[125][28] = 5'b01111; w[125][29] = 5'b01111; w[125][30] = 5'b01111; w[125][31] = 5'b00000; w[125][32] = 5'b10000; w[125][33] = 5'b10000; w[125][34] = 5'b10000; w[125][35] = 5'b10000; w[125][36] = 5'b10000; w[125][37] = 5'b10000; w[125][38] = 5'b00000; w[125][39] = 5'b01111; w[125][40] = 5'b01111; w[125][41] = 5'b01111; w[125][42] = 5'b01111; w[125][43] = 5'b01111; w[125][44] = 5'b01111; w[125][45] = 5'b10000; w[125][46] = 5'b10000; w[125][47] = 5'b10000; w[125][48] = 5'b10000; w[125][49] = 5'b10000; w[125][50] = 5'b10000; w[125][51] = 5'b10000; w[125][52] = 5'b10000; w[125][53] = 5'b01111; w[125][54] = 5'b01111; w[125][55] = 5'b01111; w[125][56] = 5'b01111; w[125][57] = 5'b01111; w[125][58] = 5'b01111; w[125][59] = 5'b00000; w[125][60] = 5'b00000; w[125][61] = 5'b01111; w[125][62] = 5'b10000; w[125][63] = 5'b00000; w[125][64] = 5'b01111; w[125][65] = 5'b00000; w[125][66] = 5'b00000; w[125][67] = 5'b01111; w[125][68] = 5'b01111; w[125][69] = 5'b01111; w[125][70] = 5'b01111; w[125][71] = 5'b01111; w[125][72] = 5'b01111; w[125][73] = 5'b00000; w[125][74] = 5'b01111; w[125][75] = 5'b01111; w[125][76] = 5'b10000; w[125][77] = 5'b00000; w[125][78] = 5'b01111; w[125][79] = 5'b01111; w[125][80] = 5'b00000; w[125][81] = 5'b01111; w[125][82] = 5'b01111; w[125][83] = 5'b01111; w[125][84] = 5'b01111; w[125][85] = 5'b01111; w[125][86] = 5'b01111; w[125][87] = 5'b00000; w[125][88] = 5'b01111; w[125][89] = 5'b01111; w[125][90] = 5'b10000; w[125][91] = 5'b10000; w[125][92] = 5'b01111; w[125][93] = 5'b01111; w[125][94] = 5'b01111; w[125][95] = 5'b01111; w[125][96] = 5'b01111; w[125][97] = 5'b01111; w[125][98] = 5'b01111; w[125][99] = 5'b01111; w[125][100] = 5'b01111; w[125][101] = 5'b00000; w[125][102] = 5'b01111; w[125][103] = 5'b01111; w[125][104] = 5'b10000; w[125][105] = 5'b10000; w[125][106] = 5'b01111; w[125][107] = 5'b00000; w[125][108] = 5'b00000; w[125][109] = 5'b01111; w[125][110] = 5'b01111; w[125][111] = 5'b01111; w[125][112] = 5'b01111; w[125][113] = 5'b01111; w[125][114] = 5'b01111; w[125][115] = 5'b00000; w[125][116] = 5'b01111; w[125][117] = 5'b01111; w[125][118] = 5'b10000; w[125][119] = 5'b10000; w[125][120] = 5'b00000; w[125][121] = 5'b00000; w[125][122] = 5'b00000; w[125][123] = 5'b01111; w[125][124] = 5'b01111; w[125][125] = 5'b00000; w[125][126] = 5'b01111; w[125][127] = 5'b01111; w[125][128] = 5'b01111; w[125][129] = 5'b00000; w[125][130] = 5'b01111; w[125][131] = 5'b01111; w[125][132] = 5'b00000; w[125][133] = 5'b10000; w[125][134] = 5'b01111; w[125][135] = 5'b01111; w[125][136] = 5'b00000; w[125][137] = 5'b01111; w[125][138] = 5'b01111; w[125][139] = 5'b01111; w[125][140] = 5'b01111; w[125][141] = 5'b01111; w[125][142] = 5'b01111; w[125][143] = 5'b00000; w[125][144] = 5'b00000; w[125][145] = 5'b01111; w[125][146] = 5'b00000; w[125][147] = 5'b10000; w[125][148] = 5'b01111; w[125][149] = 5'b00000; w[125][150] = 5'b00000; w[125][151] = 5'b01111; w[125][152] = 5'b01111; w[125][153] = 5'b01111; w[125][154] = 5'b01111; w[125][155] = 5'b01111; w[125][156] = 5'b01111; w[125][157] = 5'b00000; w[125][158] = 5'b00000; w[125][159] = 5'b00000; w[125][160] = 5'b10000; w[125][161] = 5'b10000; w[125][162] = 5'b10000; w[125][163] = 5'b00000; w[125][164] = 5'b00000; w[125][165] = 5'b01111; w[125][166] = 5'b01111; w[125][167] = 5'b01111; w[125][168] = 5'b01111; w[125][169] = 5'b01111; w[125][170] = 5'b01111; w[125][171] = 5'b01111; w[125][172] = 5'b00000; w[125][173] = 5'b00000; w[125][174] = 5'b10000; w[125][175] = 5'b10000; w[125][176] = 5'b10000; w[125][177] = 5'b00000; w[125][178] = 5'b01111; w[125][179] = 5'b01111; w[125][180] = 5'b01111; w[125][181] = 5'b01111; w[125][182] = 5'b01111; w[125][183] = 5'b01111; w[125][184] = 5'b01111; w[125][185] = 5'b01111; w[125][186] = 5'b01111; w[125][187] = 5'b01111; w[125][188] = 5'b01111; w[125][189] = 5'b01111; w[125][190] = 5'b01111; w[125][191] = 5'b01111; w[125][192] = 5'b01111; w[125][193] = 5'b01111; w[125][194] = 5'b01111; w[125][195] = 5'b01111; w[125][196] = 5'b01111; w[125][197] = 5'b01111; w[125][198] = 5'b01111; w[125][199] = 5'b01111; w[125][200] = 5'b01111; w[125][201] = 5'b01111; w[125][202] = 5'b01111; w[125][203] = 5'b01111; w[125][204] = 5'b01111; w[125][205] = 5'b01111; w[125][206] = 5'b01111; w[125][207] = 5'b01111; w[125][208] = 5'b01111; w[125][209] = 5'b01111; 
w[126][0] = 5'b01111; w[126][1] = 5'b01111; w[126][2] = 5'b01111; w[126][3] = 5'b01111; w[126][4] = 5'b01111; w[126][5] = 5'b01111; w[126][6] = 5'b01111; w[126][7] = 5'b01111; w[126][8] = 5'b01111; w[126][9] = 5'b01111; w[126][10] = 5'b01111; w[126][11] = 5'b01111; w[126][12] = 5'b01111; w[126][13] = 5'b01111; w[126][14] = 5'b01111; w[126][15] = 5'b01111; w[126][16] = 5'b01111; w[126][17] = 5'b01111; w[126][18] = 5'b01111; w[126][19] = 5'b01111; w[126][20] = 5'b01111; w[126][21] = 5'b01111; w[126][22] = 5'b01111; w[126][23] = 5'b01111; w[126][24] = 5'b01111; w[126][25] = 5'b01111; w[126][26] = 5'b01111; w[126][27] = 5'b01111; w[126][28] = 5'b01111; w[126][29] = 5'b01111; w[126][30] = 5'b01111; w[126][31] = 5'b00000; w[126][32] = 5'b10000; w[126][33] = 5'b10000; w[126][34] = 5'b10000; w[126][35] = 5'b10000; w[126][36] = 5'b10000; w[126][37] = 5'b10000; w[126][38] = 5'b00000; w[126][39] = 5'b01111; w[126][40] = 5'b01111; w[126][41] = 5'b01111; w[126][42] = 5'b01111; w[126][43] = 5'b01111; w[126][44] = 5'b01111; w[126][45] = 5'b10000; w[126][46] = 5'b10000; w[126][47] = 5'b10000; w[126][48] = 5'b10000; w[126][49] = 5'b10000; w[126][50] = 5'b10000; w[126][51] = 5'b10000; w[126][52] = 5'b10000; w[126][53] = 5'b01111; w[126][54] = 5'b01111; w[126][55] = 5'b01111; w[126][56] = 5'b01111; w[126][57] = 5'b01111; w[126][58] = 5'b01111; w[126][59] = 5'b00000; w[126][60] = 5'b00000; w[126][61] = 5'b01111; w[126][62] = 5'b10000; w[126][63] = 5'b00000; w[126][64] = 5'b01111; w[126][65] = 5'b00000; w[126][66] = 5'b00000; w[126][67] = 5'b01111; w[126][68] = 5'b01111; w[126][69] = 5'b01111; w[126][70] = 5'b01111; w[126][71] = 5'b01111; w[126][72] = 5'b01111; w[126][73] = 5'b00000; w[126][74] = 5'b01111; w[126][75] = 5'b01111; w[126][76] = 5'b10000; w[126][77] = 5'b00000; w[126][78] = 5'b01111; w[126][79] = 5'b01111; w[126][80] = 5'b00000; w[126][81] = 5'b01111; w[126][82] = 5'b01111; w[126][83] = 5'b01111; w[126][84] = 5'b01111; w[126][85] = 5'b01111; w[126][86] = 5'b01111; w[126][87] = 5'b00000; w[126][88] = 5'b01111; w[126][89] = 5'b01111; w[126][90] = 5'b10000; w[126][91] = 5'b10000; w[126][92] = 5'b01111; w[126][93] = 5'b01111; w[126][94] = 5'b01111; w[126][95] = 5'b01111; w[126][96] = 5'b01111; w[126][97] = 5'b01111; w[126][98] = 5'b01111; w[126][99] = 5'b01111; w[126][100] = 5'b01111; w[126][101] = 5'b00000; w[126][102] = 5'b01111; w[126][103] = 5'b01111; w[126][104] = 5'b10000; w[126][105] = 5'b10000; w[126][106] = 5'b01111; w[126][107] = 5'b00000; w[126][108] = 5'b00000; w[126][109] = 5'b01111; w[126][110] = 5'b01111; w[126][111] = 5'b01111; w[126][112] = 5'b01111; w[126][113] = 5'b01111; w[126][114] = 5'b01111; w[126][115] = 5'b00000; w[126][116] = 5'b01111; w[126][117] = 5'b01111; w[126][118] = 5'b10000; w[126][119] = 5'b10000; w[126][120] = 5'b00000; w[126][121] = 5'b00000; w[126][122] = 5'b00000; w[126][123] = 5'b01111; w[126][124] = 5'b01111; w[126][125] = 5'b01111; w[126][126] = 5'b00000; w[126][127] = 5'b01111; w[126][128] = 5'b01111; w[126][129] = 5'b00000; w[126][130] = 5'b01111; w[126][131] = 5'b01111; w[126][132] = 5'b00000; w[126][133] = 5'b10000; w[126][134] = 5'b01111; w[126][135] = 5'b01111; w[126][136] = 5'b00000; w[126][137] = 5'b01111; w[126][138] = 5'b01111; w[126][139] = 5'b01111; w[126][140] = 5'b01111; w[126][141] = 5'b01111; w[126][142] = 5'b01111; w[126][143] = 5'b00000; w[126][144] = 5'b00000; w[126][145] = 5'b01111; w[126][146] = 5'b00000; w[126][147] = 5'b10000; w[126][148] = 5'b01111; w[126][149] = 5'b00000; w[126][150] = 5'b00000; w[126][151] = 5'b01111; w[126][152] = 5'b01111; w[126][153] = 5'b01111; w[126][154] = 5'b01111; w[126][155] = 5'b01111; w[126][156] = 5'b01111; w[126][157] = 5'b00000; w[126][158] = 5'b00000; w[126][159] = 5'b00000; w[126][160] = 5'b10000; w[126][161] = 5'b10000; w[126][162] = 5'b10000; w[126][163] = 5'b00000; w[126][164] = 5'b00000; w[126][165] = 5'b01111; w[126][166] = 5'b01111; w[126][167] = 5'b01111; w[126][168] = 5'b01111; w[126][169] = 5'b01111; w[126][170] = 5'b01111; w[126][171] = 5'b01111; w[126][172] = 5'b00000; w[126][173] = 5'b00000; w[126][174] = 5'b10000; w[126][175] = 5'b10000; w[126][176] = 5'b10000; w[126][177] = 5'b00000; w[126][178] = 5'b01111; w[126][179] = 5'b01111; w[126][180] = 5'b01111; w[126][181] = 5'b01111; w[126][182] = 5'b01111; w[126][183] = 5'b01111; w[126][184] = 5'b01111; w[126][185] = 5'b01111; w[126][186] = 5'b01111; w[126][187] = 5'b01111; w[126][188] = 5'b01111; w[126][189] = 5'b01111; w[126][190] = 5'b01111; w[126][191] = 5'b01111; w[126][192] = 5'b01111; w[126][193] = 5'b01111; w[126][194] = 5'b01111; w[126][195] = 5'b01111; w[126][196] = 5'b01111; w[126][197] = 5'b01111; w[126][198] = 5'b01111; w[126][199] = 5'b01111; w[126][200] = 5'b01111; w[126][201] = 5'b01111; w[126][202] = 5'b01111; w[126][203] = 5'b01111; w[126][204] = 5'b01111; w[126][205] = 5'b01111; w[126][206] = 5'b01111; w[126][207] = 5'b01111; w[126][208] = 5'b01111; w[126][209] = 5'b01111; 
w[127][0] = 5'b01111; w[127][1] = 5'b01111; w[127][2] = 5'b01111; w[127][3] = 5'b01111; w[127][4] = 5'b01111; w[127][5] = 5'b01111; w[127][6] = 5'b01111; w[127][7] = 5'b01111; w[127][8] = 5'b01111; w[127][9] = 5'b01111; w[127][10] = 5'b01111; w[127][11] = 5'b01111; w[127][12] = 5'b01111; w[127][13] = 5'b01111; w[127][14] = 5'b01111; w[127][15] = 5'b01111; w[127][16] = 5'b01111; w[127][17] = 5'b01111; w[127][18] = 5'b01111; w[127][19] = 5'b01111; w[127][20] = 5'b01111; w[127][21] = 5'b01111; w[127][22] = 5'b01111; w[127][23] = 5'b01111; w[127][24] = 5'b01111; w[127][25] = 5'b01111; w[127][26] = 5'b01111; w[127][27] = 5'b01111; w[127][28] = 5'b01111; w[127][29] = 5'b01111; w[127][30] = 5'b01111; w[127][31] = 5'b00000; w[127][32] = 5'b10000; w[127][33] = 5'b10000; w[127][34] = 5'b10000; w[127][35] = 5'b10000; w[127][36] = 5'b10000; w[127][37] = 5'b10000; w[127][38] = 5'b00000; w[127][39] = 5'b01111; w[127][40] = 5'b01111; w[127][41] = 5'b01111; w[127][42] = 5'b01111; w[127][43] = 5'b01111; w[127][44] = 5'b01111; w[127][45] = 5'b10000; w[127][46] = 5'b10000; w[127][47] = 5'b10000; w[127][48] = 5'b10000; w[127][49] = 5'b10000; w[127][50] = 5'b10000; w[127][51] = 5'b10000; w[127][52] = 5'b10000; w[127][53] = 5'b01111; w[127][54] = 5'b01111; w[127][55] = 5'b01111; w[127][56] = 5'b01111; w[127][57] = 5'b01111; w[127][58] = 5'b01111; w[127][59] = 5'b00000; w[127][60] = 5'b00000; w[127][61] = 5'b01111; w[127][62] = 5'b10000; w[127][63] = 5'b00000; w[127][64] = 5'b01111; w[127][65] = 5'b00000; w[127][66] = 5'b00000; w[127][67] = 5'b01111; w[127][68] = 5'b01111; w[127][69] = 5'b01111; w[127][70] = 5'b01111; w[127][71] = 5'b01111; w[127][72] = 5'b01111; w[127][73] = 5'b00000; w[127][74] = 5'b01111; w[127][75] = 5'b01111; w[127][76] = 5'b10000; w[127][77] = 5'b00000; w[127][78] = 5'b01111; w[127][79] = 5'b01111; w[127][80] = 5'b00000; w[127][81] = 5'b01111; w[127][82] = 5'b01111; w[127][83] = 5'b01111; w[127][84] = 5'b01111; w[127][85] = 5'b01111; w[127][86] = 5'b01111; w[127][87] = 5'b00000; w[127][88] = 5'b01111; w[127][89] = 5'b01111; w[127][90] = 5'b10000; w[127][91] = 5'b10000; w[127][92] = 5'b01111; w[127][93] = 5'b01111; w[127][94] = 5'b01111; w[127][95] = 5'b01111; w[127][96] = 5'b01111; w[127][97] = 5'b01111; w[127][98] = 5'b01111; w[127][99] = 5'b01111; w[127][100] = 5'b01111; w[127][101] = 5'b00000; w[127][102] = 5'b01111; w[127][103] = 5'b01111; w[127][104] = 5'b10000; w[127][105] = 5'b10000; w[127][106] = 5'b01111; w[127][107] = 5'b00000; w[127][108] = 5'b00000; w[127][109] = 5'b01111; w[127][110] = 5'b01111; w[127][111] = 5'b01111; w[127][112] = 5'b01111; w[127][113] = 5'b01111; w[127][114] = 5'b01111; w[127][115] = 5'b00000; w[127][116] = 5'b01111; w[127][117] = 5'b01111; w[127][118] = 5'b10000; w[127][119] = 5'b10000; w[127][120] = 5'b00000; w[127][121] = 5'b00000; w[127][122] = 5'b00000; w[127][123] = 5'b01111; w[127][124] = 5'b01111; w[127][125] = 5'b01111; w[127][126] = 5'b01111; w[127][127] = 5'b00000; w[127][128] = 5'b01111; w[127][129] = 5'b00000; w[127][130] = 5'b01111; w[127][131] = 5'b01111; w[127][132] = 5'b00000; w[127][133] = 5'b10000; w[127][134] = 5'b01111; w[127][135] = 5'b01111; w[127][136] = 5'b00000; w[127][137] = 5'b01111; w[127][138] = 5'b01111; w[127][139] = 5'b01111; w[127][140] = 5'b01111; w[127][141] = 5'b01111; w[127][142] = 5'b01111; w[127][143] = 5'b00000; w[127][144] = 5'b00000; w[127][145] = 5'b01111; w[127][146] = 5'b00000; w[127][147] = 5'b10000; w[127][148] = 5'b01111; w[127][149] = 5'b00000; w[127][150] = 5'b00000; w[127][151] = 5'b01111; w[127][152] = 5'b01111; w[127][153] = 5'b01111; w[127][154] = 5'b01111; w[127][155] = 5'b01111; w[127][156] = 5'b01111; w[127][157] = 5'b00000; w[127][158] = 5'b00000; w[127][159] = 5'b00000; w[127][160] = 5'b10000; w[127][161] = 5'b10000; w[127][162] = 5'b10000; w[127][163] = 5'b00000; w[127][164] = 5'b00000; w[127][165] = 5'b01111; w[127][166] = 5'b01111; w[127][167] = 5'b01111; w[127][168] = 5'b01111; w[127][169] = 5'b01111; w[127][170] = 5'b01111; w[127][171] = 5'b01111; w[127][172] = 5'b00000; w[127][173] = 5'b00000; w[127][174] = 5'b10000; w[127][175] = 5'b10000; w[127][176] = 5'b10000; w[127][177] = 5'b00000; w[127][178] = 5'b01111; w[127][179] = 5'b01111; w[127][180] = 5'b01111; w[127][181] = 5'b01111; w[127][182] = 5'b01111; w[127][183] = 5'b01111; w[127][184] = 5'b01111; w[127][185] = 5'b01111; w[127][186] = 5'b01111; w[127][187] = 5'b01111; w[127][188] = 5'b01111; w[127][189] = 5'b01111; w[127][190] = 5'b01111; w[127][191] = 5'b01111; w[127][192] = 5'b01111; w[127][193] = 5'b01111; w[127][194] = 5'b01111; w[127][195] = 5'b01111; w[127][196] = 5'b01111; w[127][197] = 5'b01111; w[127][198] = 5'b01111; w[127][199] = 5'b01111; w[127][200] = 5'b01111; w[127][201] = 5'b01111; w[127][202] = 5'b01111; w[127][203] = 5'b01111; w[127][204] = 5'b01111; w[127][205] = 5'b01111; w[127][206] = 5'b01111; w[127][207] = 5'b01111; w[127][208] = 5'b01111; w[127][209] = 5'b01111; 
w[128][0] = 5'b01111; w[128][1] = 5'b01111; w[128][2] = 5'b01111; w[128][3] = 5'b01111; w[128][4] = 5'b01111; w[128][5] = 5'b01111; w[128][6] = 5'b01111; w[128][7] = 5'b01111; w[128][8] = 5'b01111; w[128][9] = 5'b01111; w[128][10] = 5'b01111; w[128][11] = 5'b01111; w[128][12] = 5'b01111; w[128][13] = 5'b01111; w[128][14] = 5'b01111; w[128][15] = 5'b01111; w[128][16] = 5'b01111; w[128][17] = 5'b01111; w[128][18] = 5'b01111; w[128][19] = 5'b01111; w[128][20] = 5'b01111; w[128][21] = 5'b01111; w[128][22] = 5'b01111; w[128][23] = 5'b01111; w[128][24] = 5'b01111; w[128][25] = 5'b01111; w[128][26] = 5'b01111; w[128][27] = 5'b01111; w[128][28] = 5'b01111; w[128][29] = 5'b01111; w[128][30] = 5'b00000; w[128][31] = 5'b10000; w[128][32] = 5'b00000; w[128][33] = 5'b10000; w[128][34] = 5'b00000; w[128][35] = 5'b00000; w[128][36] = 5'b00000; w[128][37] = 5'b00000; w[128][38] = 5'b10000; w[128][39] = 5'b00000; w[128][40] = 5'b01111; w[128][41] = 5'b01111; w[128][42] = 5'b01111; w[128][43] = 5'b01111; w[128][44] = 5'b00000; w[128][45] = 5'b00000; w[128][46] = 5'b00000; w[128][47] = 5'b10000; w[128][48] = 5'b00000; w[128][49] = 5'b00000; w[128][50] = 5'b00000; w[128][51] = 5'b00000; w[128][52] = 5'b00000; w[128][53] = 5'b00000; w[128][54] = 5'b01111; w[128][55] = 5'b01111; w[128][56] = 5'b01111; w[128][57] = 5'b01111; w[128][58] = 5'b01111; w[128][59] = 5'b01111; w[128][60] = 5'b01111; w[128][61] = 5'b00000; w[128][62] = 5'b10000; w[128][63] = 5'b10000; w[128][64] = 5'b01111; w[128][65] = 5'b01111; w[128][66] = 5'b01111; w[128][67] = 5'b01111; w[128][68] = 5'b01111; w[128][69] = 5'b01111; w[128][70] = 5'b01111; w[128][71] = 5'b01111; w[128][72] = 5'b01111; w[128][73] = 5'b01111; w[128][74] = 5'b00000; w[128][75] = 5'b00000; w[128][76] = 5'b10000; w[128][77] = 5'b10000; w[128][78] = 5'b01111; w[128][79] = 5'b00000; w[128][80] = 5'b01111; w[128][81] = 5'b01111; w[128][82] = 5'b01111; w[128][83] = 5'b01111; w[128][84] = 5'b01111; w[128][85] = 5'b01111; w[128][86] = 5'b01111; w[128][87] = 5'b01111; w[128][88] = 5'b00000; w[128][89] = 5'b00000; w[128][90] = 5'b10000; w[128][91] = 5'b10000; w[128][92] = 5'b01111; w[128][93] = 5'b00000; w[128][94] = 5'b00000; w[128][95] = 5'b01111; w[128][96] = 5'b01111; w[128][97] = 5'b01111; w[128][98] = 5'b01111; w[128][99] = 5'b01111; w[128][100] = 5'b01111; w[128][101] = 5'b01111; w[128][102] = 5'b00000; w[128][103] = 5'b01111; w[128][104] = 5'b10000; w[128][105] = 5'b10000; w[128][106] = 5'b01111; w[128][107] = 5'b01111; w[128][108] = 5'b01111; w[128][109] = 5'b01111; w[128][110] = 5'b01111; w[128][111] = 5'b01111; w[128][112] = 5'b01111; w[128][113] = 5'b01111; w[128][114] = 5'b01111; w[128][115] = 5'b01111; w[128][116] = 5'b00000; w[128][117] = 5'b01111; w[128][118] = 5'b10000; w[128][119] = 5'b10000; w[128][120] = 5'b01111; w[128][121] = 5'b01111; w[128][122] = 5'b01111; w[128][123] = 5'b01111; w[128][124] = 5'b01111; w[128][125] = 5'b01111; w[128][126] = 5'b01111; w[128][127] = 5'b01111; w[128][128] = 5'b00000; w[128][129] = 5'b01111; w[128][130] = 5'b00000; w[128][131] = 5'b01111; w[128][132] = 5'b10000; w[128][133] = 5'b10000; w[128][134] = 5'b00000; w[128][135] = 5'b00000; w[128][136] = 5'b01111; w[128][137] = 5'b01111; w[128][138] = 5'b01111; w[128][139] = 5'b01111; w[128][140] = 5'b01111; w[128][141] = 5'b01111; w[128][142] = 5'b01111; w[128][143] = 5'b01111; w[128][144] = 5'b01111; w[128][145] = 5'b01111; w[128][146] = 5'b10000; w[128][147] = 5'b10000; w[128][148] = 5'b00000; w[128][149] = 5'b01111; w[128][150] = 5'b01111; w[128][151] = 5'b01111; w[128][152] = 5'b01111; w[128][153] = 5'b01111; w[128][154] = 5'b01111; w[128][155] = 5'b01111; w[128][156] = 5'b01111; w[128][157] = 5'b01111; w[128][158] = 5'b01111; w[128][159] = 5'b01111; w[128][160] = 5'b00000; w[128][161] = 5'b00000; w[128][162] = 5'b00000; w[128][163] = 5'b01111; w[128][164] = 5'b01111; w[128][165] = 5'b01111; w[128][166] = 5'b01111; w[128][167] = 5'b01111; w[128][168] = 5'b01111; w[128][169] = 5'b01111; w[128][170] = 5'b01111; w[128][171] = 5'b00000; w[128][172] = 5'b01111; w[128][173] = 5'b01111; w[128][174] = 5'b00000; w[128][175] = 5'b00000; w[128][176] = 5'b00000; w[128][177] = 5'b01111; w[128][178] = 5'b00000; w[128][179] = 5'b01111; w[128][180] = 5'b01111; w[128][181] = 5'b01111; w[128][182] = 5'b01111; w[128][183] = 5'b01111; w[128][184] = 5'b01111; w[128][185] = 5'b01111; w[128][186] = 5'b01111; w[128][187] = 5'b01111; w[128][188] = 5'b01111; w[128][189] = 5'b01111; w[128][190] = 5'b01111; w[128][191] = 5'b01111; w[128][192] = 5'b01111; w[128][193] = 5'b01111; w[128][194] = 5'b01111; w[128][195] = 5'b01111; w[128][196] = 5'b01111; w[128][197] = 5'b01111; w[128][198] = 5'b01111; w[128][199] = 5'b01111; w[128][200] = 5'b01111; w[128][201] = 5'b01111; w[128][202] = 5'b01111; w[128][203] = 5'b01111; w[128][204] = 5'b01111; w[128][205] = 5'b01111; w[128][206] = 5'b01111; w[128][207] = 5'b01111; w[128][208] = 5'b01111; w[128][209] = 5'b01111; 
w[129][0] = 5'b00000; w[129][1] = 5'b00000; w[129][2] = 5'b00000; w[129][3] = 5'b00000; w[129][4] = 5'b00000; w[129][5] = 5'b00000; w[129][6] = 5'b00000; w[129][7] = 5'b00000; w[129][8] = 5'b00000; w[129][9] = 5'b00000; w[129][10] = 5'b00000; w[129][11] = 5'b00000; w[129][12] = 5'b00000; w[129][13] = 5'b00000; w[129][14] = 5'b00000; w[129][15] = 5'b00000; w[129][16] = 5'b00000; w[129][17] = 5'b00000; w[129][18] = 5'b00000; w[129][19] = 5'b00000; w[129][20] = 5'b00000; w[129][21] = 5'b00000; w[129][22] = 5'b00000; w[129][23] = 5'b00000; w[129][24] = 5'b00000; w[129][25] = 5'b00000; w[129][26] = 5'b00000; w[129][27] = 5'b00000; w[129][28] = 5'b00000; w[129][29] = 5'b00000; w[129][30] = 5'b10000; w[129][31] = 5'b00000; w[129][32] = 5'b01111; w[129][33] = 5'b00000; w[129][34] = 5'b10000; w[129][35] = 5'b10000; w[129][36] = 5'b10000; w[129][37] = 5'b01111; w[129][38] = 5'b00000; w[129][39] = 5'b10000; w[129][40] = 5'b00000; w[129][41] = 5'b00000; w[129][42] = 5'b00000; w[129][43] = 5'b00000; w[129][44] = 5'b10000; w[129][45] = 5'b01111; w[129][46] = 5'b01111; w[129][47] = 5'b00000; w[129][48] = 5'b10000; w[129][49] = 5'b10000; w[129][50] = 5'b10000; w[129][51] = 5'b01111; w[129][52] = 5'b01111; w[129][53] = 5'b10000; w[129][54] = 5'b00000; w[129][55] = 5'b00000; w[129][56] = 5'b00000; w[129][57] = 5'b00000; w[129][58] = 5'b01111; w[129][59] = 5'b01111; w[129][60] = 5'b01111; w[129][61] = 5'b01111; w[129][62] = 5'b10000; w[129][63] = 5'b10000; w[129][64] = 5'b00000; w[129][65] = 5'b01111; w[129][66] = 5'b01111; w[129][67] = 5'b01111; w[129][68] = 5'b00000; w[129][69] = 5'b00000; w[129][70] = 5'b00000; w[129][71] = 5'b00000; w[129][72] = 5'b01111; w[129][73] = 5'b01111; w[129][74] = 5'b01111; w[129][75] = 5'b01111; w[129][76] = 5'b10000; w[129][77] = 5'b10000; w[129][78] = 5'b00000; w[129][79] = 5'b01111; w[129][80] = 5'b01111; w[129][81] = 5'b01111; w[129][82] = 5'b00000; w[129][83] = 5'b00000; w[129][84] = 5'b00000; w[129][85] = 5'b00000; w[129][86] = 5'b01111; w[129][87] = 5'b01111; w[129][88] = 5'b01111; w[129][89] = 5'b01111; w[129][90] = 5'b10000; w[129][91] = 5'b10000; w[129][92] = 5'b00000; w[129][93] = 5'b01111; w[129][94] = 5'b01111; w[129][95] = 5'b00000; w[129][96] = 5'b00000; w[129][97] = 5'b00000; w[129][98] = 5'b00000; w[129][99] = 5'b00000; w[129][100] = 5'b01111; w[129][101] = 5'b01111; w[129][102] = 5'b01111; w[129][103] = 5'b00000; w[129][104] = 5'b10000; w[129][105] = 5'b10000; w[129][106] = 5'b01111; w[129][107] = 5'b01111; w[129][108] = 5'b01111; w[129][109] = 5'b01111; w[129][110] = 5'b00000; w[129][111] = 5'b00000; w[129][112] = 5'b00000; w[129][113] = 5'b00000; w[129][114] = 5'b01111; w[129][115] = 5'b01111; w[129][116] = 5'b01111; w[129][117] = 5'b00000; w[129][118] = 5'b10000; w[129][119] = 5'b10000; w[129][120] = 5'b01111; w[129][121] = 5'b01111; w[129][122] = 5'b01111; w[129][123] = 5'b01111; w[129][124] = 5'b00000; w[129][125] = 5'b00000; w[129][126] = 5'b00000; w[129][127] = 5'b00000; w[129][128] = 5'b01111; w[129][129] = 5'b00000; w[129][130] = 5'b01111; w[129][131] = 5'b00000; w[129][132] = 5'b10000; w[129][133] = 5'b10000; w[129][134] = 5'b01111; w[129][135] = 5'b01111; w[129][136] = 5'b01111; w[129][137] = 5'b01111; w[129][138] = 5'b00000; w[129][139] = 5'b00000; w[129][140] = 5'b00000; w[129][141] = 5'b00000; w[129][142] = 5'b01111; w[129][143] = 5'b01111; w[129][144] = 5'b01111; w[129][145] = 5'b00000; w[129][146] = 5'b10000; w[129][147] = 5'b10000; w[129][148] = 5'b01111; w[129][149] = 5'b01111; w[129][150] = 5'b01111; w[129][151] = 5'b01111; w[129][152] = 5'b00000; w[129][153] = 5'b00000; w[129][154] = 5'b00000; w[129][155] = 5'b00000; w[129][156] = 5'b00000; w[129][157] = 5'b01111; w[129][158] = 5'b01111; w[129][159] = 5'b00000; w[129][160] = 5'b10000; w[129][161] = 5'b10000; w[129][162] = 5'b01111; w[129][163] = 5'b01111; w[129][164] = 5'b01111; w[129][165] = 5'b00000; w[129][166] = 5'b00000; w[129][167] = 5'b00000; w[129][168] = 5'b00000; w[129][169] = 5'b00000; w[129][170] = 5'b00000; w[129][171] = 5'b01111; w[129][172] = 5'b01111; w[129][173] = 5'b00000; w[129][174] = 5'b10000; w[129][175] = 5'b10000; w[129][176] = 5'b01111; w[129][177] = 5'b01111; w[129][178] = 5'b01111; w[129][179] = 5'b00000; w[129][180] = 5'b00000; w[129][181] = 5'b00000; w[129][182] = 5'b00000; w[129][183] = 5'b00000; w[129][184] = 5'b00000; w[129][185] = 5'b00000; w[129][186] = 5'b00000; w[129][187] = 5'b00000; w[129][188] = 5'b00000; w[129][189] = 5'b00000; w[129][190] = 5'b00000; w[129][191] = 5'b00000; w[129][192] = 5'b00000; w[129][193] = 5'b00000; w[129][194] = 5'b00000; w[129][195] = 5'b00000; w[129][196] = 5'b00000; w[129][197] = 5'b00000; w[129][198] = 5'b00000; w[129][199] = 5'b00000; w[129][200] = 5'b00000; w[129][201] = 5'b00000; w[129][202] = 5'b00000; w[129][203] = 5'b00000; w[129][204] = 5'b00000; w[129][205] = 5'b00000; w[129][206] = 5'b00000; w[129][207] = 5'b00000; w[129][208] = 5'b00000; w[129][209] = 5'b00000; 
w[130][0] = 5'b01111; w[130][1] = 5'b01111; w[130][2] = 5'b01111; w[130][3] = 5'b01111; w[130][4] = 5'b01111; w[130][5] = 5'b01111; w[130][6] = 5'b01111; w[130][7] = 5'b01111; w[130][8] = 5'b01111; w[130][9] = 5'b01111; w[130][10] = 5'b01111; w[130][11] = 5'b01111; w[130][12] = 5'b01111; w[130][13] = 5'b01111; w[130][14] = 5'b01111; w[130][15] = 5'b01111; w[130][16] = 5'b01111; w[130][17] = 5'b01111; w[130][18] = 5'b01111; w[130][19] = 5'b01111; w[130][20] = 5'b01111; w[130][21] = 5'b01111; w[130][22] = 5'b01111; w[130][23] = 5'b01111; w[130][24] = 5'b01111; w[130][25] = 5'b01111; w[130][26] = 5'b01111; w[130][27] = 5'b01111; w[130][28] = 5'b01111; w[130][29] = 5'b01111; w[130][30] = 5'b00000; w[130][31] = 5'b01111; w[130][32] = 5'b00000; w[130][33] = 5'b10000; w[130][34] = 5'b10000; w[130][35] = 5'b10000; w[130][36] = 5'b10000; w[130][37] = 5'b00000; w[130][38] = 5'b01111; w[130][39] = 5'b00000; w[130][40] = 5'b01111; w[130][41] = 5'b01111; w[130][42] = 5'b01111; w[130][43] = 5'b01111; w[130][44] = 5'b00000; w[130][45] = 5'b00000; w[130][46] = 5'b00000; w[130][47] = 5'b10000; w[130][48] = 5'b10000; w[130][49] = 5'b10000; w[130][50] = 5'b10000; w[130][51] = 5'b00000; w[130][52] = 5'b00000; w[130][53] = 5'b00000; w[130][54] = 5'b01111; w[130][55] = 5'b01111; w[130][56] = 5'b01111; w[130][57] = 5'b01111; w[130][58] = 5'b00000; w[130][59] = 5'b01111; w[130][60] = 5'b01111; w[130][61] = 5'b01111; w[130][62] = 5'b00000; w[130][63] = 5'b10000; w[130][64] = 5'b01111; w[130][65] = 5'b01111; w[130][66] = 5'b01111; w[130][67] = 5'b00000; w[130][68] = 5'b01111; w[130][69] = 5'b01111; w[130][70] = 5'b01111; w[130][71] = 5'b01111; w[130][72] = 5'b00000; w[130][73] = 5'b01111; w[130][74] = 5'b01111; w[130][75] = 5'b01111; w[130][76] = 5'b00000; w[130][77] = 5'b10000; w[130][78] = 5'b01111; w[130][79] = 5'b01111; w[130][80] = 5'b01111; w[130][81] = 5'b00000; w[130][82] = 5'b01111; w[130][83] = 5'b01111; w[130][84] = 5'b01111; w[130][85] = 5'b01111; w[130][86] = 5'b00000; w[130][87] = 5'b01111; w[130][88] = 5'b01111; w[130][89] = 5'b01111; w[130][90] = 5'b00000; w[130][91] = 5'b00000; w[130][92] = 5'b01111; w[130][93] = 5'b01111; w[130][94] = 5'b01111; w[130][95] = 5'b01111; w[130][96] = 5'b01111; w[130][97] = 5'b01111; w[130][98] = 5'b01111; w[130][99] = 5'b01111; w[130][100] = 5'b00000; w[130][101] = 5'b01111; w[130][102] = 5'b01111; w[130][103] = 5'b01111; w[130][104] = 5'b00000; w[130][105] = 5'b00000; w[130][106] = 5'b00000; w[130][107] = 5'b01111; w[130][108] = 5'b01111; w[130][109] = 5'b00000; w[130][110] = 5'b01111; w[130][111] = 5'b01111; w[130][112] = 5'b01111; w[130][113] = 5'b01111; w[130][114] = 5'b00000; w[130][115] = 5'b01111; w[130][116] = 5'b01111; w[130][117] = 5'b01111; w[130][118] = 5'b00000; w[130][119] = 5'b00000; w[130][120] = 5'b01111; w[130][121] = 5'b01111; w[130][122] = 5'b01111; w[130][123] = 5'b00000; w[130][124] = 5'b01111; w[130][125] = 5'b01111; w[130][126] = 5'b01111; w[130][127] = 5'b01111; w[130][128] = 5'b00000; w[130][129] = 5'b01111; w[130][130] = 5'b00000; w[130][131] = 5'b01111; w[130][132] = 5'b10000; w[130][133] = 5'b00000; w[130][134] = 5'b01111; w[130][135] = 5'b01111; w[130][136] = 5'b01111; w[130][137] = 5'b00000; w[130][138] = 5'b01111; w[130][139] = 5'b01111; w[130][140] = 5'b01111; w[130][141] = 5'b01111; w[130][142] = 5'b00000; w[130][143] = 5'b01111; w[130][144] = 5'b01111; w[130][145] = 5'b01111; w[130][146] = 5'b10000; w[130][147] = 5'b00000; w[130][148] = 5'b01111; w[130][149] = 5'b01111; w[130][150] = 5'b01111; w[130][151] = 5'b00000; w[130][152] = 5'b01111; w[130][153] = 5'b01111; w[130][154] = 5'b01111; w[130][155] = 5'b01111; w[130][156] = 5'b01111; w[130][157] = 5'b01111; w[130][158] = 5'b01111; w[130][159] = 5'b10000; w[130][160] = 5'b10000; w[130][161] = 5'b10000; w[130][162] = 5'b00000; w[130][163] = 5'b01111; w[130][164] = 5'b01111; w[130][165] = 5'b01111; w[130][166] = 5'b01111; w[130][167] = 5'b01111; w[130][168] = 5'b01111; w[130][169] = 5'b01111; w[130][170] = 5'b01111; w[130][171] = 5'b01111; w[130][172] = 5'b01111; w[130][173] = 5'b10000; w[130][174] = 5'b10000; w[130][175] = 5'b10000; w[130][176] = 5'b00000; w[130][177] = 5'b01111; w[130][178] = 5'b01111; w[130][179] = 5'b01111; w[130][180] = 5'b01111; w[130][181] = 5'b01111; w[130][182] = 5'b01111; w[130][183] = 5'b01111; w[130][184] = 5'b01111; w[130][185] = 5'b01111; w[130][186] = 5'b01111; w[130][187] = 5'b01111; w[130][188] = 5'b01111; w[130][189] = 5'b01111; w[130][190] = 5'b01111; w[130][191] = 5'b01111; w[130][192] = 5'b01111; w[130][193] = 5'b01111; w[130][194] = 5'b01111; w[130][195] = 5'b01111; w[130][196] = 5'b01111; w[130][197] = 5'b01111; w[130][198] = 5'b01111; w[130][199] = 5'b01111; w[130][200] = 5'b01111; w[130][201] = 5'b01111; w[130][202] = 5'b01111; w[130][203] = 5'b01111; w[130][204] = 5'b01111; w[130][205] = 5'b01111; w[130][206] = 5'b01111; w[130][207] = 5'b01111; w[130][208] = 5'b01111; w[130][209] = 5'b01111; 
w[131][0] = 5'b01111; w[131][1] = 5'b01111; w[131][2] = 5'b01111; w[131][3] = 5'b01111; w[131][4] = 5'b01111; w[131][5] = 5'b01111; w[131][6] = 5'b01111; w[131][7] = 5'b01111; w[131][8] = 5'b01111; w[131][9] = 5'b01111; w[131][10] = 5'b01111; w[131][11] = 5'b01111; w[131][12] = 5'b01111; w[131][13] = 5'b01111; w[131][14] = 5'b01111; w[131][15] = 5'b01111; w[131][16] = 5'b01111; w[131][17] = 5'b01111; w[131][18] = 5'b01111; w[131][19] = 5'b01111; w[131][20] = 5'b01111; w[131][21] = 5'b01111; w[131][22] = 5'b01111; w[131][23] = 5'b01111; w[131][24] = 5'b01111; w[131][25] = 5'b01111; w[131][26] = 5'b01111; w[131][27] = 5'b01111; w[131][28] = 5'b01111; w[131][29] = 5'b01111; w[131][30] = 5'b01111; w[131][31] = 5'b00000; w[131][32] = 5'b10000; w[131][33] = 5'b10000; w[131][34] = 5'b10000; w[131][35] = 5'b10000; w[131][36] = 5'b10000; w[131][37] = 5'b10000; w[131][38] = 5'b00000; w[131][39] = 5'b01111; w[131][40] = 5'b01111; w[131][41] = 5'b01111; w[131][42] = 5'b01111; w[131][43] = 5'b01111; w[131][44] = 5'b01111; w[131][45] = 5'b10000; w[131][46] = 5'b10000; w[131][47] = 5'b10000; w[131][48] = 5'b10000; w[131][49] = 5'b10000; w[131][50] = 5'b10000; w[131][51] = 5'b10000; w[131][52] = 5'b10000; w[131][53] = 5'b01111; w[131][54] = 5'b01111; w[131][55] = 5'b01111; w[131][56] = 5'b01111; w[131][57] = 5'b01111; w[131][58] = 5'b01111; w[131][59] = 5'b00000; w[131][60] = 5'b00000; w[131][61] = 5'b01111; w[131][62] = 5'b10000; w[131][63] = 5'b00000; w[131][64] = 5'b01111; w[131][65] = 5'b00000; w[131][66] = 5'b00000; w[131][67] = 5'b01111; w[131][68] = 5'b01111; w[131][69] = 5'b01111; w[131][70] = 5'b01111; w[131][71] = 5'b01111; w[131][72] = 5'b01111; w[131][73] = 5'b00000; w[131][74] = 5'b01111; w[131][75] = 5'b01111; w[131][76] = 5'b10000; w[131][77] = 5'b00000; w[131][78] = 5'b01111; w[131][79] = 5'b01111; w[131][80] = 5'b00000; w[131][81] = 5'b01111; w[131][82] = 5'b01111; w[131][83] = 5'b01111; w[131][84] = 5'b01111; w[131][85] = 5'b01111; w[131][86] = 5'b01111; w[131][87] = 5'b00000; w[131][88] = 5'b01111; w[131][89] = 5'b01111; w[131][90] = 5'b10000; w[131][91] = 5'b10000; w[131][92] = 5'b01111; w[131][93] = 5'b01111; w[131][94] = 5'b01111; w[131][95] = 5'b01111; w[131][96] = 5'b01111; w[131][97] = 5'b01111; w[131][98] = 5'b01111; w[131][99] = 5'b01111; w[131][100] = 5'b01111; w[131][101] = 5'b00000; w[131][102] = 5'b01111; w[131][103] = 5'b01111; w[131][104] = 5'b10000; w[131][105] = 5'b10000; w[131][106] = 5'b01111; w[131][107] = 5'b00000; w[131][108] = 5'b00000; w[131][109] = 5'b01111; w[131][110] = 5'b01111; w[131][111] = 5'b01111; w[131][112] = 5'b01111; w[131][113] = 5'b01111; w[131][114] = 5'b01111; w[131][115] = 5'b00000; w[131][116] = 5'b01111; w[131][117] = 5'b01111; w[131][118] = 5'b10000; w[131][119] = 5'b10000; w[131][120] = 5'b00000; w[131][121] = 5'b00000; w[131][122] = 5'b00000; w[131][123] = 5'b01111; w[131][124] = 5'b01111; w[131][125] = 5'b01111; w[131][126] = 5'b01111; w[131][127] = 5'b01111; w[131][128] = 5'b01111; w[131][129] = 5'b00000; w[131][130] = 5'b01111; w[131][131] = 5'b00000; w[131][132] = 5'b00000; w[131][133] = 5'b10000; w[131][134] = 5'b01111; w[131][135] = 5'b01111; w[131][136] = 5'b00000; w[131][137] = 5'b01111; w[131][138] = 5'b01111; w[131][139] = 5'b01111; w[131][140] = 5'b01111; w[131][141] = 5'b01111; w[131][142] = 5'b01111; w[131][143] = 5'b00000; w[131][144] = 5'b00000; w[131][145] = 5'b01111; w[131][146] = 5'b00000; w[131][147] = 5'b10000; w[131][148] = 5'b01111; w[131][149] = 5'b00000; w[131][150] = 5'b00000; w[131][151] = 5'b01111; w[131][152] = 5'b01111; w[131][153] = 5'b01111; w[131][154] = 5'b01111; w[131][155] = 5'b01111; w[131][156] = 5'b01111; w[131][157] = 5'b00000; w[131][158] = 5'b00000; w[131][159] = 5'b00000; w[131][160] = 5'b10000; w[131][161] = 5'b10000; w[131][162] = 5'b10000; w[131][163] = 5'b00000; w[131][164] = 5'b00000; w[131][165] = 5'b01111; w[131][166] = 5'b01111; w[131][167] = 5'b01111; w[131][168] = 5'b01111; w[131][169] = 5'b01111; w[131][170] = 5'b01111; w[131][171] = 5'b01111; w[131][172] = 5'b00000; w[131][173] = 5'b00000; w[131][174] = 5'b10000; w[131][175] = 5'b10000; w[131][176] = 5'b10000; w[131][177] = 5'b00000; w[131][178] = 5'b01111; w[131][179] = 5'b01111; w[131][180] = 5'b01111; w[131][181] = 5'b01111; w[131][182] = 5'b01111; w[131][183] = 5'b01111; w[131][184] = 5'b01111; w[131][185] = 5'b01111; w[131][186] = 5'b01111; w[131][187] = 5'b01111; w[131][188] = 5'b01111; w[131][189] = 5'b01111; w[131][190] = 5'b01111; w[131][191] = 5'b01111; w[131][192] = 5'b01111; w[131][193] = 5'b01111; w[131][194] = 5'b01111; w[131][195] = 5'b01111; w[131][196] = 5'b01111; w[131][197] = 5'b01111; w[131][198] = 5'b01111; w[131][199] = 5'b01111; w[131][200] = 5'b01111; w[131][201] = 5'b01111; w[131][202] = 5'b01111; w[131][203] = 5'b01111; w[131][204] = 5'b01111; w[131][205] = 5'b01111; w[131][206] = 5'b01111; w[131][207] = 5'b01111; w[131][208] = 5'b01111; w[131][209] = 5'b01111; 
w[132][0] = 5'b00000; w[132][1] = 5'b00000; w[132][2] = 5'b00000; w[132][3] = 5'b00000; w[132][4] = 5'b00000; w[132][5] = 5'b00000; w[132][6] = 5'b00000; w[132][7] = 5'b00000; w[132][8] = 5'b00000; w[132][9] = 5'b00000; w[132][10] = 5'b00000; w[132][11] = 5'b00000; w[132][12] = 5'b00000; w[132][13] = 5'b00000; w[132][14] = 5'b00000; w[132][15] = 5'b00000; w[132][16] = 5'b00000; w[132][17] = 5'b00000; w[132][18] = 5'b00000; w[132][19] = 5'b00000; w[132][20] = 5'b00000; w[132][21] = 5'b00000; w[132][22] = 5'b00000; w[132][23] = 5'b00000; w[132][24] = 5'b00000; w[132][25] = 5'b00000; w[132][26] = 5'b00000; w[132][27] = 5'b00000; w[132][28] = 5'b00000; w[132][29] = 5'b00000; w[132][30] = 5'b01111; w[132][31] = 5'b00000; w[132][32] = 5'b10000; w[132][33] = 5'b00000; w[132][34] = 5'b01111; w[132][35] = 5'b01111; w[132][36] = 5'b01111; w[132][37] = 5'b10000; w[132][38] = 5'b00000; w[132][39] = 5'b01111; w[132][40] = 5'b00000; w[132][41] = 5'b00000; w[132][42] = 5'b00000; w[132][43] = 5'b00000; w[132][44] = 5'b01111; w[132][45] = 5'b10000; w[132][46] = 5'b10000; w[132][47] = 5'b00000; w[132][48] = 5'b01111; w[132][49] = 5'b01111; w[132][50] = 5'b01111; w[132][51] = 5'b10000; w[132][52] = 5'b10000; w[132][53] = 5'b01111; w[132][54] = 5'b00000; w[132][55] = 5'b00000; w[132][56] = 5'b00000; w[132][57] = 5'b00000; w[132][58] = 5'b10000; w[132][59] = 5'b10000; w[132][60] = 5'b10000; w[132][61] = 5'b10000; w[132][62] = 5'b01111; w[132][63] = 5'b01111; w[132][64] = 5'b00000; w[132][65] = 5'b10000; w[132][66] = 5'b10000; w[132][67] = 5'b10000; w[132][68] = 5'b00000; w[132][69] = 5'b00000; w[132][70] = 5'b00000; w[132][71] = 5'b00000; w[132][72] = 5'b10000; w[132][73] = 5'b10000; w[132][74] = 5'b10000; w[132][75] = 5'b10000; w[132][76] = 5'b01111; w[132][77] = 5'b01111; w[132][78] = 5'b00000; w[132][79] = 5'b10000; w[132][80] = 5'b10000; w[132][81] = 5'b10000; w[132][82] = 5'b00000; w[132][83] = 5'b00000; w[132][84] = 5'b00000; w[132][85] = 5'b00000; w[132][86] = 5'b10000; w[132][87] = 5'b10000; w[132][88] = 5'b10000; w[132][89] = 5'b10000; w[132][90] = 5'b01111; w[132][91] = 5'b01111; w[132][92] = 5'b00000; w[132][93] = 5'b10000; w[132][94] = 5'b10000; w[132][95] = 5'b00000; w[132][96] = 5'b00000; w[132][97] = 5'b00000; w[132][98] = 5'b00000; w[132][99] = 5'b00000; w[132][100] = 5'b10000; w[132][101] = 5'b10000; w[132][102] = 5'b10000; w[132][103] = 5'b00000; w[132][104] = 5'b01111; w[132][105] = 5'b01111; w[132][106] = 5'b10000; w[132][107] = 5'b10000; w[132][108] = 5'b10000; w[132][109] = 5'b10000; w[132][110] = 5'b00000; w[132][111] = 5'b00000; w[132][112] = 5'b00000; w[132][113] = 5'b00000; w[132][114] = 5'b10000; w[132][115] = 5'b10000; w[132][116] = 5'b10000; w[132][117] = 5'b00000; w[132][118] = 5'b01111; w[132][119] = 5'b01111; w[132][120] = 5'b10000; w[132][121] = 5'b10000; w[132][122] = 5'b10000; w[132][123] = 5'b10000; w[132][124] = 5'b00000; w[132][125] = 5'b00000; w[132][126] = 5'b00000; w[132][127] = 5'b00000; w[132][128] = 5'b10000; w[132][129] = 5'b10000; w[132][130] = 5'b10000; w[132][131] = 5'b00000; w[132][132] = 5'b00000; w[132][133] = 5'b01111; w[132][134] = 5'b10000; w[132][135] = 5'b10000; w[132][136] = 5'b10000; w[132][137] = 5'b10000; w[132][138] = 5'b00000; w[132][139] = 5'b00000; w[132][140] = 5'b00000; w[132][141] = 5'b00000; w[132][142] = 5'b10000; w[132][143] = 5'b10000; w[132][144] = 5'b10000; w[132][145] = 5'b00000; w[132][146] = 5'b01111; w[132][147] = 5'b01111; w[132][148] = 5'b10000; w[132][149] = 5'b10000; w[132][150] = 5'b10000; w[132][151] = 5'b10000; w[132][152] = 5'b00000; w[132][153] = 5'b00000; w[132][154] = 5'b00000; w[132][155] = 5'b00000; w[132][156] = 5'b00000; w[132][157] = 5'b10000; w[132][158] = 5'b10000; w[132][159] = 5'b00000; w[132][160] = 5'b01111; w[132][161] = 5'b01111; w[132][162] = 5'b10000; w[132][163] = 5'b10000; w[132][164] = 5'b10000; w[132][165] = 5'b00000; w[132][166] = 5'b00000; w[132][167] = 5'b00000; w[132][168] = 5'b00000; w[132][169] = 5'b00000; w[132][170] = 5'b00000; w[132][171] = 5'b10000; w[132][172] = 5'b10000; w[132][173] = 5'b00000; w[132][174] = 5'b01111; w[132][175] = 5'b01111; w[132][176] = 5'b10000; w[132][177] = 5'b10000; w[132][178] = 5'b10000; w[132][179] = 5'b00000; w[132][180] = 5'b00000; w[132][181] = 5'b00000; w[132][182] = 5'b00000; w[132][183] = 5'b00000; w[132][184] = 5'b00000; w[132][185] = 5'b00000; w[132][186] = 5'b00000; w[132][187] = 5'b00000; w[132][188] = 5'b00000; w[132][189] = 5'b00000; w[132][190] = 5'b00000; w[132][191] = 5'b00000; w[132][192] = 5'b00000; w[132][193] = 5'b00000; w[132][194] = 5'b00000; w[132][195] = 5'b00000; w[132][196] = 5'b00000; w[132][197] = 5'b00000; w[132][198] = 5'b00000; w[132][199] = 5'b00000; w[132][200] = 5'b00000; w[132][201] = 5'b00000; w[132][202] = 5'b00000; w[132][203] = 5'b00000; w[132][204] = 5'b00000; w[132][205] = 5'b00000; w[132][206] = 5'b00000; w[132][207] = 5'b00000; w[132][208] = 5'b00000; w[132][209] = 5'b00000; 
w[133][0] = 5'b10000; w[133][1] = 5'b10000; w[133][2] = 5'b10000; w[133][3] = 5'b10000; w[133][4] = 5'b10000; w[133][5] = 5'b10000; w[133][6] = 5'b10000; w[133][7] = 5'b10000; w[133][8] = 5'b10000; w[133][9] = 5'b10000; w[133][10] = 5'b10000; w[133][11] = 5'b10000; w[133][12] = 5'b10000; w[133][13] = 5'b10000; w[133][14] = 5'b10000; w[133][15] = 5'b10000; w[133][16] = 5'b10000; w[133][17] = 5'b10000; w[133][18] = 5'b10000; w[133][19] = 5'b10000; w[133][20] = 5'b10000; w[133][21] = 5'b10000; w[133][22] = 5'b10000; w[133][23] = 5'b10000; w[133][24] = 5'b10000; w[133][25] = 5'b10000; w[133][26] = 5'b10000; w[133][27] = 5'b10000; w[133][28] = 5'b10000; w[133][29] = 5'b10000; w[133][30] = 5'b00000; w[133][31] = 5'b01111; w[133][32] = 5'b00000; w[133][33] = 5'b01111; w[133][34] = 5'b00000; w[133][35] = 5'b00000; w[133][36] = 5'b00000; w[133][37] = 5'b00000; w[133][38] = 5'b01111; w[133][39] = 5'b00000; w[133][40] = 5'b10000; w[133][41] = 5'b10000; w[133][42] = 5'b10000; w[133][43] = 5'b10000; w[133][44] = 5'b00000; w[133][45] = 5'b00000; w[133][46] = 5'b00000; w[133][47] = 5'b01111; w[133][48] = 5'b00000; w[133][49] = 5'b00000; w[133][50] = 5'b00000; w[133][51] = 5'b00000; w[133][52] = 5'b00000; w[133][53] = 5'b00000; w[133][54] = 5'b10000; w[133][55] = 5'b10000; w[133][56] = 5'b10000; w[133][57] = 5'b10000; w[133][58] = 5'b10000; w[133][59] = 5'b10000; w[133][60] = 5'b10000; w[133][61] = 5'b00000; w[133][62] = 5'b01111; w[133][63] = 5'b01111; w[133][64] = 5'b10000; w[133][65] = 5'b10000; w[133][66] = 5'b10000; w[133][67] = 5'b10000; w[133][68] = 5'b10000; w[133][69] = 5'b10000; w[133][70] = 5'b10000; w[133][71] = 5'b10000; w[133][72] = 5'b10000; w[133][73] = 5'b10000; w[133][74] = 5'b00000; w[133][75] = 5'b00000; w[133][76] = 5'b01111; w[133][77] = 5'b01111; w[133][78] = 5'b10000; w[133][79] = 5'b00000; w[133][80] = 5'b10000; w[133][81] = 5'b10000; w[133][82] = 5'b10000; w[133][83] = 5'b10000; w[133][84] = 5'b10000; w[133][85] = 5'b10000; w[133][86] = 5'b10000; w[133][87] = 5'b10000; w[133][88] = 5'b00000; w[133][89] = 5'b00000; w[133][90] = 5'b01111; w[133][91] = 5'b01111; w[133][92] = 5'b10000; w[133][93] = 5'b00000; w[133][94] = 5'b00000; w[133][95] = 5'b10000; w[133][96] = 5'b10000; w[133][97] = 5'b10000; w[133][98] = 5'b10000; w[133][99] = 5'b10000; w[133][100] = 5'b10000; w[133][101] = 5'b10000; w[133][102] = 5'b00000; w[133][103] = 5'b10000; w[133][104] = 5'b01111; w[133][105] = 5'b01111; w[133][106] = 5'b10000; w[133][107] = 5'b10000; w[133][108] = 5'b10000; w[133][109] = 5'b10000; w[133][110] = 5'b10000; w[133][111] = 5'b10000; w[133][112] = 5'b10000; w[133][113] = 5'b10000; w[133][114] = 5'b10000; w[133][115] = 5'b10000; w[133][116] = 5'b00000; w[133][117] = 5'b10000; w[133][118] = 5'b01111; w[133][119] = 5'b01111; w[133][120] = 5'b10000; w[133][121] = 5'b10000; w[133][122] = 5'b10000; w[133][123] = 5'b10000; w[133][124] = 5'b10000; w[133][125] = 5'b10000; w[133][126] = 5'b10000; w[133][127] = 5'b10000; w[133][128] = 5'b10000; w[133][129] = 5'b10000; w[133][130] = 5'b00000; w[133][131] = 5'b10000; w[133][132] = 5'b01111; w[133][133] = 5'b00000; w[133][134] = 5'b00000; w[133][135] = 5'b00000; w[133][136] = 5'b10000; w[133][137] = 5'b10000; w[133][138] = 5'b10000; w[133][139] = 5'b10000; w[133][140] = 5'b10000; w[133][141] = 5'b10000; w[133][142] = 5'b10000; w[133][143] = 5'b10000; w[133][144] = 5'b10000; w[133][145] = 5'b10000; w[133][146] = 5'b01111; w[133][147] = 5'b01111; w[133][148] = 5'b00000; w[133][149] = 5'b10000; w[133][150] = 5'b10000; w[133][151] = 5'b10000; w[133][152] = 5'b10000; w[133][153] = 5'b10000; w[133][154] = 5'b10000; w[133][155] = 5'b10000; w[133][156] = 5'b10000; w[133][157] = 5'b10000; w[133][158] = 5'b10000; w[133][159] = 5'b10000; w[133][160] = 5'b00000; w[133][161] = 5'b00000; w[133][162] = 5'b00000; w[133][163] = 5'b10000; w[133][164] = 5'b10000; w[133][165] = 5'b10000; w[133][166] = 5'b10000; w[133][167] = 5'b10000; w[133][168] = 5'b10000; w[133][169] = 5'b10000; w[133][170] = 5'b10000; w[133][171] = 5'b00000; w[133][172] = 5'b10000; w[133][173] = 5'b10000; w[133][174] = 5'b00000; w[133][175] = 5'b00000; w[133][176] = 5'b00000; w[133][177] = 5'b10000; w[133][178] = 5'b00000; w[133][179] = 5'b10000; w[133][180] = 5'b10000; w[133][181] = 5'b10000; w[133][182] = 5'b10000; w[133][183] = 5'b10000; w[133][184] = 5'b10000; w[133][185] = 5'b10000; w[133][186] = 5'b10000; w[133][187] = 5'b10000; w[133][188] = 5'b10000; w[133][189] = 5'b10000; w[133][190] = 5'b10000; w[133][191] = 5'b10000; w[133][192] = 5'b10000; w[133][193] = 5'b10000; w[133][194] = 5'b10000; w[133][195] = 5'b10000; w[133][196] = 5'b10000; w[133][197] = 5'b10000; w[133][198] = 5'b10000; w[133][199] = 5'b10000; w[133][200] = 5'b10000; w[133][201] = 5'b10000; w[133][202] = 5'b10000; w[133][203] = 5'b10000; w[133][204] = 5'b10000; w[133][205] = 5'b10000; w[133][206] = 5'b10000; w[133][207] = 5'b10000; w[133][208] = 5'b10000; w[133][209] = 5'b10000; 
w[134][0] = 5'b01111; w[134][1] = 5'b01111; w[134][2] = 5'b01111; w[134][3] = 5'b01111; w[134][4] = 5'b01111; w[134][5] = 5'b01111; w[134][6] = 5'b01111; w[134][7] = 5'b01111; w[134][8] = 5'b01111; w[134][9] = 5'b01111; w[134][10] = 5'b01111; w[134][11] = 5'b01111; w[134][12] = 5'b01111; w[134][13] = 5'b01111; w[134][14] = 5'b01111; w[134][15] = 5'b01111; w[134][16] = 5'b01111; w[134][17] = 5'b01111; w[134][18] = 5'b01111; w[134][19] = 5'b01111; w[134][20] = 5'b01111; w[134][21] = 5'b01111; w[134][22] = 5'b01111; w[134][23] = 5'b01111; w[134][24] = 5'b01111; w[134][25] = 5'b01111; w[134][26] = 5'b01111; w[134][27] = 5'b01111; w[134][28] = 5'b01111; w[134][29] = 5'b01111; w[134][30] = 5'b00000; w[134][31] = 5'b01111; w[134][32] = 5'b00000; w[134][33] = 5'b10000; w[134][34] = 5'b10000; w[134][35] = 5'b10000; w[134][36] = 5'b10000; w[134][37] = 5'b00000; w[134][38] = 5'b01111; w[134][39] = 5'b00000; w[134][40] = 5'b01111; w[134][41] = 5'b01111; w[134][42] = 5'b01111; w[134][43] = 5'b01111; w[134][44] = 5'b00000; w[134][45] = 5'b00000; w[134][46] = 5'b00000; w[134][47] = 5'b10000; w[134][48] = 5'b10000; w[134][49] = 5'b10000; w[134][50] = 5'b10000; w[134][51] = 5'b00000; w[134][52] = 5'b00000; w[134][53] = 5'b00000; w[134][54] = 5'b01111; w[134][55] = 5'b01111; w[134][56] = 5'b01111; w[134][57] = 5'b01111; w[134][58] = 5'b00000; w[134][59] = 5'b01111; w[134][60] = 5'b01111; w[134][61] = 5'b01111; w[134][62] = 5'b00000; w[134][63] = 5'b10000; w[134][64] = 5'b01111; w[134][65] = 5'b01111; w[134][66] = 5'b01111; w[134][67] = 5'b00000; w[134][68] = 5'b01111; w[134][69] = 5'b01111; w[134][70] = 5'b01111; w[134][71] = 5'b01111; w[134][72] = 5'b00000; w[134][73] = 5'b01111; w[134][74] = 5'b01111; w[134][75] = 5'b01111; w[134][76] = 5'b00000; w[134][77] = 5'b10000; w[134][78] = 5'b01111; w[134][79] = 5'b01111; w[134][80] = 5'b01111; w[134][81] = 5'b00000; w[134][82] = 5'b01111; w[134][83] = 5'b01111; w[134][84] = 5'b01111; w[134][85] = 5'b01111; w[134][86] = 5'b00000; w[134][87] = 5'b01111; w[134][88] = 5'b01111; w[134][89] = 5'b01111; w[134][90] = 5'b00000; w[134][91] = 5'b00000; w[134][92] = 5'b01111; w[134][93] = 5'b01111; w[134][94] = 5'b01111; w[134][95] = 5'b01111; w[134][96] = 5'b01111; w[134][97] = 5'b01111; w[134][98] = 5'b01111; w[134][99] = 5'b01111; w[134][100] = 5'b00000; w[134][101] = 5'b01111; w[134][102] = 5'b01111; w[134][103] = 5'b01111; w[134][104] = 5'b00000; w[134][105] = 5'b00000; w[134][106] = 5'b00000; w[134][107] = 5'b01111; w[134][108] = 5'b01111; w[134][109] = 5'b00000; w[134][110] = 5'b01111; w[134][111] = 5'b01111; w[134][112] = 5'b01111; w[134][113] = 5'b01111; w[134][114] = 5'b00000; w[134][115] = 5'b01111; w[134][116] = 5'b01111; w[134][117] = 5'b01111; w[134][118] = 5'b00000; w[134][119] = 5'b00000; w[134][120] = 5'b01111; w[134][121] = 5'b01111; w[134][122] = 5'b01111; w[134][123] = 5'b00000; w[134][124] = 5'b01111; w[134][125] = 5'b01111; w[134][126] = 5'b01111; w[134][127] = 5'b01111; w[134][128] = 5'b00000; w[134][129] = 5'b01111; w[134][130] = 5'b01111; w[134][131] = 5'b01111; w[134][132] = 5'b10000; w[134][133] = 5'b00000; w[134][134] = 5'b00000; w[134][135] = 5'b01111; w[134][136] = 5'b01111; w[134][137] = 5'b00000; w[134][138] = 5'b01111; w[134][139] = 5'b01111; w[134][140] = 5'b01111; w[134][141] = 5'b01111; w[134][142] = 5'b00000; w[134][143] = 5'b01111; w[134][144] = 5'b01111; w[134][145] = 5'b01111; w[134][146] = 5'b10000; w[134][147] = 5'b00000; w[134][148] = 5'b01111; w[134][149] = 5'b01111; w[134][150] = 5'b01111; w[134][151] = 5'b00000; w[134][152] = 5'b01111; w[134][153] = 5'b01111; w[134][154] = 5'b01111; w[134][155] = 5'b01111; w[134][156] = 5'b01111; w[134][157] = 5'b01111; w[134][158] = 5'b01111; w[134][159] = 5'b10000; w[134][160] = 5'b10000; w[134][161] = 5'b10000; w[134][162] = 5'b00000; w[134][163] = 5'b01111; w[134][164] = 5'b01111; w[134][165] = 5'b01111; w[134][166] = 5'b01111; w[134][167] = 5'b01111; w[134][168] = 5'b01111; w[134][169] = 5'b01111; w[134][170] = 5'b01111; w[134][171] = 5'b01111; w[134][172] = 5'b01111; w[134][173] = 5'b10000; w[134][174] = 5'b10000; w[134][175] = 5'b10000; w[134][176] = 5'b00000; w[134][177] = 5'b01111; w[134][178] = 5'b01111; w[134][179] = 5'b01111; w[134][180] = 5'b01111; w[134][181] = 5'b01111; w[134][182] = 5'b01111; w[134][183] = 5'b01111; w[134][184] = 5'b01111; w[134][185] = 5'b01111; w[134][186] = 5'b01111; w[134][187] = 5'b01111; w[134][188] = 5'b01111; w[134][189] = 5'b01111; w[134][190] = 5'b01111; w[134][191] = 5'b01111; w[134][192] = 5'b01111; w[134][193] = 5'b01111; w[134][194] = 5'b01111; w[134][195] = 5'b01111; w[134][196] = 5'b01111; w[134][197] = 5'b01111; w[134][198] = 5'b01111; w[134][199] = 5'b01111; w[134][200] = 5'b01111; w[134][201] = 5'b01111; w[134][202] = 5'b01111; w[134][203] = 5'b01111; w[134][204] = 5'b01111; w[134][205] = 5'b01111; w[134][206] = 5'b01111; w[134][207] = 5'b01111; w[134][208] = 5'b01111; w[134][209] = 5'b01111; 
w[135][0] = 5'b01111; w[135][1] = 5'b01111; w[135][2] = 5'b01111; w[135][3] = 5'b01111; w[135][4] = 5'b01111; w[135][5] = 5'b01111; w[135][6] = 5'b01111; w[135][7] = 5'b01111; w[135][8] = 5'b01111; w[135][9] = 5'b01111; w[135][10] = 5'b01111; w[135][11] = 5'b01111; w[135][12] = 5'b01111; w[135][13] = 5'b01111; w[135][14] = 5'b01111; w[135][15] = 5'b01111; w[135][16] = 5'b01111; w[135][17] = 5'b01111; w[135][18] = 5'b01111; w[135][19] = 5'b01111; w[135][20] = 5'b01111; w[135][21] = 5'b01111; w[135][22] = 5'b01111; w[135][23] = 5'b01111; w[135][24] = 5'b01111; w[135][25] = 5'b01111; w[135][26] = 5'b01111; w[135][27] = 5'b01111; w[135][28] = 5'b01111; w[135][29] = 5'b01111; w[135][30] = 5'b00000; w[135][31] = 5'b01111; w[135][32] = 5'b00000; w[135][33] = 5'b10000; w[135][34] = 5'b10000; w[135][35] = 5'b10000; w[135][36] = 5'b10000; w[135][37] = 5'b00000; w[135][38] = 5'b01111; w[135][39] = 5'b00000; w[135][40] = 5'b01111; w[135][41] = 5'b01111; w[135][42] = 5'b01111; w[135][43] = 5'b01111; w[135][44] = 5'b00000; w[135][45] = 5'b00000; w[135][46] = 5'b00000; w[135][47] = 5'b10000; w[135][48] = 5'b10000; w[135][49] = 5'b10000; w[135][50] = 5'b10000; w[135][51] = 5'b00000; w[135][52] = 5'b00000; w[135][53] = 5'b00000; w[135][54] = 5'b01111; w[135][55] = 5'b01111; w[135][56] = 5'b01111; w[135][57] = 5'b01111; w[135][58] = 5'b00000; w[135][59] = 5'b01111; w[135][60] = 5'b01111; w[135][61] = 5'b01111; w[135][62] = 5'b00000; w[135][63] = 5'b10000; w[135][64] = 5'b01111; w[135][65] = 5'b01111; w[135][66] = 5'b01111; w[135][67] = 5'b00000; w[135][68] = 5'b01111; w[135][69] = 5'b01111; w[135][70] = 5'b01111; w[135][71] = 5'b01111; w[135][72] = 5'b00000; w[135][73] = 5'b01111; w[135][74] = 5'b01111; w[135][75] = 5'b01111; w[135][76] = 5'b00000; w[135][77] = 5'b10000; w[135][78] = 5'b01111; w[135][79] = 5'b01111; w[135][80] = 5'b01111; w[135][81] = 5'b00000; w[135][82] = 5'b01111; w[135][83] = 5'b01111; w[135][84] = 5'b01111; w[135][85] = 5'b01111; w[135][86] = 5'b00000; w[135][87] = 5'b01111; w[135][88] = 5'b01111; w[135][89] = 5'b01111; w[135][90] = 5'b00000; w[135][91] = 5'b00000; w[135][92] = 5'b01111; w[135][93] = 5'b01111; w[135][94] = 5'b01111; w[135][95] = 5'b01111; w[135][96] = 5'b01111; w[135][97] = 5'b01111; w[135][98] = 5'b01111; w[135][99] = 5'b01111; w[135][100] = 5'b00000; w[135][101] = 5'b01111; w[135][102] = 5'b01111; w[135][103] = 5'b01111; w[135][104] = 5'b00000; w[135][105] = 5'b00000; w[135][106] = 5'b00000; w[135][107] = 5'b01111; w[135][108] = 5'b01111; w[135][109] = 5'b00000; w[135][110] = 5'b01111; w[135][111] = 5'b01111; w[135][112] = 5'b01111; w[135][113] = 5'b01111; w[135][114] = 5'b00000; w[135][115] = 5'b01111; w[135][116] = 5'b01111; w[135][117] = 5'b01111; w[135][118] = 5'b00000; w[135][119] = 5'b00000; w[135][120] = 5'b01111; w[135][121] = 5'b01111; w[135][122] = 5'b01111; w[135][123] = 5'b00000; w[135][124] = 5'b01111; w[135][125] = 5'b01111; w[135][126] = 5'b01111; w[135][127] = 5'b01111; w[135][128] = 5'b00000; w[135][129] = 5'b01111; w[135][130] = 5'b01111; w[135][131] = 5'b01111; w[135][132] = 5'b10000; w[135][133] = 5'b00000; w[135][134] = 5'b01111; w[135][135] = 5'b00000; w[135][136] = 5'b01111; w[135][137] = 5'b00000; w[135][138] = 5'b01111; w[135][139] = 5'b01111; w[135][140] = 5'b01111; w[135][141] = 5'b01111; w[135][142] = 5'b00000; w[135][143] = 5'b01111; w[135][144] = 5'b01111; w[135][145] = 5'b01111; w[135][146] = 5'b10000; w[135][147] = 5'b00000; w[135][148] = 5'b01111; w[135][149] = 5'b01111; w[135][150] = 5'b01111; w[135][151] = 5'b00000; w[135][152] = 5'b01111; w[135][153] = 5'b01111; w[135][154] = 5'b01111; w[135][155] = 5'b01111; w[135][156] = 5'b01111; w[135][157] = 5'b01111; w[135][158] = 5'b01111; w[135][159] = 5'b10000; w[135][160] = 5'b10000; w[135][161] = 5'b10000; w[135][162] = 5'b00000; w[135][163] = 5'b01111; w[135][164] = 5'b01111; w[135][165] = 5'b01111; w[135][166] = 5'b01111; w[135][167] = 5'b01111; w[135][168] = 5'b01111; w[135][169] = 5'b01111; w[135][170] = 5'b01111; w[135][171] = 5'b01111; w[135][172] = 5'b01111; w[135][173] = 5'b10000; w[135][174] = 5'b10000; w[135][175] = 5'b10000; w[135][176] = 5'b00000; w[135][177] = 5'b01111; w[135][178] = 5'b01111; w[135][179] = 5'b01111; w[135][180] = 5'b01111; w[135][181] = 5'b01111; w[135][182] = 5'b01111; w[135][183] = 5'b01111; w[135][184] = 5'b01111; w[135][185] = 5'b01111; w[135][186] = 5'b01111; w[135][187] = 5'b01111; w[135][188] = 5'b01111; w[135][189] = 5'b01111; w[135][190] = 5'b01111; w[135][191] = 5'b01111; w[135][192] = 5'b01111; w[135][193] = 5'b01111; w[135][194] = 5'b01111; w[135][195] = 5'b01111; w[135][196] = 5'b01111; w[135][197] = 5'b01111; w[135][198] = 5'b01111; w[135][199] = 5'b01111; w[135][200] = 5'b01111; w[135][201] = 5'b01111; w[135][202] = 5'b01111; w[135][203] = 5'b01111; w[135][204] = 5'b01111; w[135][205] = 5'b01111; w[135][206] = 5'b01111; w[135][207] = 5'b01111; w[135][208] = 5'b01111; w[135][209] = 5'b01111; 
w[136][0] = 5'b00000; w[136][1] = 5'b00000; w[136][2] = 5'b00000; w[136][3] = 5'b00000; w[136][4] = 5'b00000; w[136][5] = 5'b00000; w[136][6] = 5'b00000; w[136][7] = 5'b00000; w[136][8] = 5'b00000; w[136][9] = 5'b00000; w[136][10] = 5'b00000; w[136][11] = 5'b00000; w[136][12] = 5'b00000; w[136][13] = 5'b00000; w[136][14] = 5'b00000; w[136][15] = 5'b00000; w[136][16] = 5'b00000; w[136][17] = 5'b00000; w[136][18] = 5'b00000; w[136][19] = 5'b00000; w[136][20] = 5'b00000; w[136][21] = 5'b00000; w[136][22] = 5'b00000; w[136][23] = 5'b00000; w[136][24] = 5'b00000; w[136][25] = 5'b00000; w[136][26] = 5'b00000; w[136][27] = 5'b00000; w[136][28] = 5'b00000; w[136][29] = 5'b00000; w[136][30] = 5'b10000; w[136][31] = 5'b00000; w[136][32] = 5'b01111; w[136][33] = 5'b00000; w[136][34] = 5'b10000; w[136][35] = 5'b10000; w[136][36] = 5'b10000; w[136][37] = 5'b01111; w[136][38] = 5'b00000; w[136][39] = 5'b10000; w[136][40] = 5'b00000; w[136][41] = 5'b00000; w[136][42] = 5'b00000; w[136][43] = 5'b00000; w[136][44] = 5'b10000; w[136][45] = 5'b01111; w[136][46] = 5'b01111; w[136][47] = 5'b00000; w[136][48] = 5'b10000; w[136][49] = 5'b10000; w[136][50] = 5'b10000; w[136][51] = 5'b01111; w[136][52] = 5'b01111; w[136][53] = 5'b10000; w[136][54] = 5'b00000; w[136][55] = 5'b00000; w[136][56] = 5'b00000; w[136][57] = 5'b00000; w[136][58] = 5'b01111; w[136][59] = 5'b01111; w[136][60] = 5'b01111; w[136][61] = 5'b01111; w[136][62] = 5'b10000; w[136][63] = 5'b10000; w[136][64] = 5'b00000; w[136][65] = 5'b01111; w[136][66] = 5'b01111; w[136][67] = 5'b01111; w[136][68] = 5'b00000; w[136][69] = 5'b00000; w[136][70] = 5'b00000; w[136][71] = 5'b00000; w[136][72] = 5'b01111; w[136][73] = 5'b01111; w[136][74] = 5'b01111; w[136][75] = 5'b01111; w[136][76] = 5'b10000; w[136][77] = 5'b10000; w[136][78] = 5'b00000; w[136][79] = 5'b01111; w[136][80] = 5'b01111; w[136][81] = 5'b01111; w[136][82] = 5'b00000; w[136][83] = 5'b00000; w[136][84] = 5'b00000; w[136][85] = 5'b00000; w[136][86] = 5'b01111; w[136][87] = 5'b01111; w[136][88] = 5'b01111; w[136][89] = 5'b01111; w[136][90] = 5'b10000; w[136][91] = 5'b10000; w[136][92] = 5'b00000; w[136][93] = 5'b01111; w[136][94] = 5'b01111; w[136][95] = 5'b00000; w[136][96] = 5'b00000; w[136][97] = 5'b00000; w[136][98] = 5'b00000; w[136][99] = 5'b00000; w[136][100] = 5'b01111; w[136][101] = 5'b01111; w[136][102] = 5'b01111; w[136][103] = 5'b00000; w[136][104] = 5'b10000; w[136][105] = 5'b10000; w[136][106] = 5'b01111; w[136][107] = 5'b01111; w[136][108] = 5'b01111; w[136][109] = 5'b01111; w[136][110] = 5'b00000; w[136][111] = 5'b00000; w[136][112] = 5'b00000; w[136][113] = 5'b00000; w[136][114] = 5'b01111; w[136][115] = 5'b01111; w[136][116] = 5'b01111; w[136][117] = 5'b00000; w[136][118] = 5'b10000; w[136][119] = 5'b10000; w[136][120] = 5'b01111; w[136][121] = 5'b01111; w[136][122] = 5'b01111; w[136][123] = 5'b01111; w[136][124] = 5'b00000; w[136][125] = 5'b00000; w[136][126] = 5'b00000; w[136][127] = 5'b00000; w[136][128] = 5'b01111; w[136][129] = 5'b01111; w[136][130] = 5'b01111; w[136][131] = 5'b00000; w[136][132] = 5'b10000; w[136][133] = 5'b10000; w[136][134] = 5'b01111; w[136][135] = 5'b01111; w[136][136] = 5'b00000; w[136][137] = 5'b01111; w[136][138] = 5'b00000; w[136][139] = 5'b00000; w[136][140] = 5'b00000; w[136][141] = 5'b00000; w[136][142] = 5'b01111; w[136][143] = 5'b01111; w[136][144] = 5'b01111; w[136][145] = 5'b00000; w[136][146] = 5'b10000; w[136][147] = 5'b10000; w[136][148] = 5'b01111; w[136][149] = 5'b01111; w[136][150] = 5'b01111; w[136][151] = 5'b01111; w[136][152] = 5'b00000; w[136][153] = 5'b00000; w[136][154] = 5'b00000; w[136][155] = 5'b00000; w[136][156] = 5'b00000; w[136][157] = 5'b01111; w[136][158] = 5'b01111; w[136][159] = 5'b00000; w[136][160] = 5'b10000; w[136][161] = 5'b10000; w[136][162] = 5'b01111; w[136][163] = 5'b01111; w[136][164] = 5'b01111; w[136][165] = 5'b00000; w[136][166] = 5'b00000; w[136][167] = 5'b00000; w[136][168] = 5'b00000; w[136][169] = 5'b00000; w[136][170] = 5'b00000; w[136][171] = 5'b01111; w[136][172] = 5'b01111; w[136][173] = 5'b00000; w[136][174] = 5'b10000; w[136][175] = 5'b10000; w[136][176] = 5'b01111; w[136][177] = 5'b01111; w[136][178] = 5'b01111; w[136][179] = 5'b00000; w[136][180] = 5'b00000; w[136][181] = 5'b00000; w[136][182] = 5'b00000; w[136][183] = 5'b00000; w[136][184] = 5'b00000; w[136][185] = 5'b00000; w[136][186] = 5'b00000; w[136][187] = 5'b00000; w[136][188] = 5'b00000; w[136][189] = 5'b00000; w[136][190] = 5'b00000; w[136][191] = 5'b00000; w[136][192] = 5'b00000; w[136][193] = 5'b00000; w[136][194] = 5'b00000; w[136][195] = 5'b00000; w[136][196] = 5'b00000; w[136][197] = 5'b00000; w[136][198] = 5'b00000; w[136][199] = 5'b00000; w[136][200] = 5'b00000; w[136][201] = 5'b00000; w[136][202] = 5'b00000; w[136][203] = 5'b00000; w[136][204] = 5'b00000; w[136][205] = 5'b00000; w[136][206] = 5'b00000; w[136][207] = 5'b00000; w[136][208] = 5'b00000; w[136][209] = 5'b00000; 
w[137][0] = 5'b01111; w[137][1] = 5'b01111; w[137][2] = 5'b01111; w[137][3] = 5'b01111; w[137][4] = 5'b01111; w[137][5] = 5'b01111; w[137][6] = 5'b01111; w[137][7] = 5'b01111; w[137][8] = 5'b01111; w[137][9] = 5'b01111; w[137][10] = 5'b01111; w[137][11] = 5'b01111; w[137][12] = 5'b01111; w[137][13] = 5'b01111; w[137][14] = 5'b01111; w[137][15] = 5'b01111; w[137][16] = 5'b01111; w[137][17] = 5'b01111; w[137][18] = 5'b01111; w[137][19] = 5'b01111; w[137][20] = 5'b01111; w[137][21] = 5'b01111; w[137][22] = 5'b01111; w[137][23] = 5'b01111; w[137][24] = 5'b01111; w[137][25] = 5'b01111; w[137][26] = 5'b01111; w[137][27] = 5'b01111; w[137][28] = 5'b01111; w[137][29] = 5'b01111; w[137][30] = 5'b00000; w[137][31] = 5'b10000; w[137][32] = 5'b00000; w[137][33] = 5'b10000; w[137][34] = 5'b00000; w[137][35] = 5'b00000; w[137][36] = 5'b00000; w[137][37] = 5'b00000; w[137][38] = 5'b10000; w[137][39] = 5'b00000; w[137][40] = 5'b01111; w[137][41] = 5'b01111; w[137][42] = 5'b01111; w[137][43] = 5'b01111; w[137][44] = 5'b00000; w[137][45] = 5'b00000; w[137][46] = 5'b00000; w[137][47] = 5'b10000; w[137][48] = 5'b00000; w[137][49] = 5'b00000; w[137][50] = 5'b00000; w[137][51] = 5'b00000; w[137][52] = 5'b00000; w[137][53] = 5'b00000; w[137][54] = 5'b01111; w[137][55] = 5'b01111; w[137][56] = 5'b01111; w[137][57] = 5'b01111; w[137][58] = 5'b01111; w[137][59] = 5'b01111; w[137][60] = 5'b01111; w[137][61] = 5'b00000; w[137][62] = 5'b10000; w[137][63] = 5'b10000; w[137][64] = 5'b01111; w[137][65] = 5'b01111; w[137][66] = 5'b01111; w[137][67] = 5'b01111; w[137][68] = 5'b01111; w[137][69] = 5'b01111; w[137][70] = 5'b01111; w[137][71] = 5'b01111; w[137][72] = 5'b01111; w[137][73] = 5'b01111; w[137][74] = 5'b00000; w[137][75] = 5'b00000; w[137][76] = 5'b10000; w[137][77] = 5'b10000; w[137][78] = 5'b01111; w[137][79] = 5'b00000; w[137][80] = 5'b01111; w[137][81] = 5'b01111; w[137][82] = 5'b01111; w[137][83] = 5'b01111; w[137][84] = 5'b01111; w[137][85] = 5'b01111; w[137][86] = 5'b01111; w[137][87] = 5'b01111; w[137][88] = 5'b00000; w[137][89] = 5'b00000; w[137][90] = 5'b10000; w[137][91] = 5'b10000; w[137][92] = 5'b01111; w[137][93] = 5'b00000; w[137][94] = 5'b00000; w[137][95] = 5'b01111; w[137][96] = 5'b01111; w[137][97] = 5'b01111; w[137][98] = 5'b01111; w[137][99] = 5'b01111; w[137][100] = 5'b01111; w[137][101] = 5'b01111; w[137][102] = 5'b00000; w[137][103] = 5'b01111; w[137][104] = 5'b10000; w[137][105] = 5'b10000; w[137][106] = 5'b01111; w[137][107] = 5'b01111; w[137][108] = 5'b01111; w[137][109] = 5'b01111; w[137][110] = 5'b01111; w[137][111] = 5'b01111; w[137][112] = 5'b01111; w[137][113] = 5'b01111; w[137][114] = 5'b01111; w[137][115] = 5'b01111; w[137][116] = 5'b00000; w[137][117] = 5'b01111; w[137][118] = 5'b10000; w[137][119] = 5'b10000; w[137][120] = 5'b01111; w[137][121] = 5'b01111; w[137][122] = 5'b01111; w[137][123] = 5'b01111; w[137][124] = 5'b01111; w[137][125] = 5'b01111; w[137][126] = 5'b01111; w[137][127] = 5'b01111; w[137][128] = 5'b01111; w[137][129] = 5'b01111; w[137][130] = 5'b00000; w[137][131] = 5'b01111; w[137][132] = 5'b10000; w[137][133] = 5'b10000; w[137][134] = 5'b00000; w[137][135] = 5'b00000; w[137][136] = 5'b01111; w[137][137] = 5'b00000; w[137][138] = 5'b01111; w[137][139] = 5'b01111; w[137][140] = 5'b01111; w[137][141] = 5'b01111; w[137][142] = 5'b01111; w[137][143] = 5'b01111; w[137][144] = 5'b01111; w[137][145] = 5'b01111; w[137][146] = 5'b10000; w[137][147] = 5'b10000; w[137][148] = 5'b00000; w[137][149] = 5'b01111; w[137][150] = 5'b01111; w[137][151] = 5'b01111; w[137][152] = 5'b01111; w[137][153] = 5'b01111; w[137][154] = 5'b01111; w[137][155] = 5'b01111; w[137][156] = 5'b01111; w[137][157] = 5'b01111; w[137][158] = 5'b01111; w[137][159] = 5'b01111; w[137][160] = 5'b00000; w[137][161] = 5'b00000; w[137][162] = 5'b00000; w[137][163] = 5'b01111; w[137][164] = 5'b01111; w[137][165] = 5'b01111; w[137][166] = 5'b01111; w[137][167] = 5'b01111; w[137][168] = 5'b01111; w[137][169] = 5'b01111; w[137][170] = 5'b01111; w[137][171] = 5'b00000; w[137][172] = 5'b01111; w[137][173] = 5'b01111; w[137][174] = 5'b00000; w[137][175] = 5'b00000; w[137][176] = 5'b00000; w[137][177] = 5'b01111; w[137][178] = 5'b00000; w[137][179] = 5'b01111; w[137][180] = 5'b01111; w[137][181] = 5'b01111; w[137][182] = 5'b01111; w[137][183] = 5'b01111; w[137][184] = 5'b01111; w[137][185] = 5'b01111; w[137][186] = 5'b01111; w[137][187] = 5'b01111; w[137][188] = 5'b01111; w[137][189] = 5'b01111; w[137][190] = 5'b01111; w[137][191] = 5'b01111; w[137][192] = 5'b01111; w[137][193] = 5'b01111; w[137][194] = 5'b01111; w[137][195] = 5'b01111; w[137][196] = 5'b01111; w[137][197] = 5'b01111; w[137][198] = 5'b01111; w[137][199] = 5'b01111; w[137][200] = 5'b01111; w[137][201] = 5'b01111; w[137][202] = 5'b01111; w[137][203] = 5'b01111; w[137][204] = 5'b01111; w[137][205] = 5'b01111; w[137][206] = 5'b01111; w[137][207] = 5'b01111; w[137][208] = 5'b01111; w[137][209] = 5'b01111; 
w[138][0] = 5'b01111; w[138][1] = 5'b01111; w[138][2] = 5'b01111; w[138][3] = 5'b01111; w[138][4] = 5'b01111; w[138][5] = 5'b01111; w[138][6] = 5'b01111; w[138][7] = 5'b01111; w[138][8] = 5'b01111; w[138][9] = 5'b01111; w[138][10] = 5'b01111; w[138][11] = 5'b01111; w[138][12] = 5'b01111; w[138][13] = 5'b01111; w[138][14] = 5'b01111; w[138][15] = 5'b01111; w[138][16] = 5'b01111; w[138][17] = 5'b01111; w[138][18] = 5'b01111; w[138][19] = 5'b01111; w[138][20] = 5'b01111; w[138][21] = 5'b01111; w[138][22] = 5'b01111; w[138][23] = 5'b01111; w[138][24] = 5'b01111; w[138][25] = 5'b01111; w[138][26] = 5'b01111; w[138][27] = 5'b01111; w[138][28] = 5'b01111; w[138][29] = 5'b01111; w[138][30] = 5'b01111; w[138][31] = 5'b00000; w[138][32] = 5'b10000; w[138][33] = 5'b10000; w[138][34] = 5'b10000; w[138][35] = 5'b10000; w[138][36] = 5'b10000; w[138][37] = 5'b10000; w[138][38] = 5'b00000; w[138][39] = 5'b01111; w[138][40] = 5'b01111; w[138][41] = 5'b01111; w[138][42] = 5'b01111; w[138][43] = 5'b01111; w[138][44] = 5'b01111; w[138][45] = 5'b10000; w[138][46] = 5'b10000; w[138][47] = 5'b10000; w[138][48] = 5'b10000; w[138][49] = 5'b10000; w[138][50] = 5'b10000; w[138][51] = 5'b10000; w[138][52] = 5'b10000; w[138][53] = 5'b01111; w[138][54] = 5'b01111; w[138][55] = 5'b01111; w[138][56] = 5'b01111; w[138][57] = 5'b01111; w[138][58] = 5'b01111; w[138][59] = 5'b00000; w[138][60] = 5'b00000; w[138][61] = 5'b01111; w[138][62] = 5'b10000; w[138][63] = 5'b00000; w[138][64] = 5'b01111; w[138][65] = 5'b00000; w[138][66] = 5'b00000; w[138][67] = 5'b01111; w[138][68] = 5'b01111; w[138][69] = 5'b01111; w[138][70] = 5'b01111; w[138][71] = 5'b01111; w[138][72] = 5'b01111; w[138][73] = 5'b00000; w[138][74] = 5'b01111; w[138][75] = 5'b01111; w[138][76] = 5'b10000; w[138][77] = 5'b00000; w[138][78] = 5'b01111; w[138][79] = 5'b01111; w[138][80] = 5'b00000; w[138][81] = 5'b01111; w[138][82] = 5'b01111; w[138][83] = 5'b01111; w[138][84] = 5'b01111; w[138][85] = 5'b01111; w[138][86] = 5'b01111; w[138][87] = 5'b00000; w[138][88] = 5'b01111; w[138][89] = 5'b01111; w[138][90] = 5'b10000; w[138][91] = 5'b10000; w[138][92] = 5'b01111; w[138][93] = 5'b01111; w[138][94] = 5'b01111; w[138][95] = 5'b01111; w[138][96] = 5'b01111; w[138][97] = 5'b01111; w[138][98] = 5'b01111; w[138][99] = 5'b01111; w[138][100] = 5'b01111; w[138][101] = 5'b00000; w[138][102] = 5'b01111; w[138][103] = 5'b01111; w[138][104] = 5'b10000; w[138][105] = 5'b10000; w[138][106] = 5'b01111; w[138][107] = 5'b00000; w[138][108] = 5'b00000; w[138][109] = 5'b01111; w[138][110] = 5'b01111; w[138][111] = 5'b01111; w[138][112] = 5'b01111; w[138][113] = 5'b01111; w[138][114] = 5'b01111; w[138][115] = 5'b00000; w[138][116] = 5'b01111; w[138][117] = 5'b01111; w[138][118] = 5'b10000; w[138][119] = 5'b10000; w[138][120] = 5'b00000; w[138][121] = 5'b00000; w[138][122] = 5'b00000; w[138][123] = 5'b01111; w[138][124] = 5'b01111; w[138][125] = 5'b01111; w[138][126] = 5'b01111; w[138][127] = 5'b01111; w[138][128] = 5'b01111; w[138][129] = 5'b00000; w[138][130] = 5'b01111; w[138][131] = 5'b01111; w[138][132] = 5'b00000; w[138][133] = 5'b10000; w[138][134] = 5'b01111; w[138][135] = 5'b01111; w[138][136] = 5'b00000; w[138][137] = 5'b01111; w[138][138] = 5'b00000; w[138][139] = 5'b01111; w[138][140] = 5'b01111; w[138][141] = 5'b01111; w[138][142] = 5'b01111; w[138][143] = 5'b00000; w[138][144] = 5'b00000; w[138][145] = 5'b01111; w[138][146] = 5'b00000; w[138][147] = 5'b10000; w[138][148] = 5'b01111; w[138][149] = 5'b00000; w[138][150] = 5'b00000; w[138][151] = 5'b01111; w[138][152] = 5'b01111; w[138][153] = 5'b01111; w[138][154] = 5'b01111; w[138][155] = 5'b01111; w[138][156] = 5'b01111; w[138][157] = 5'b00000; w[138][158] = 5'b00000; w[138][159] = 5'b00000; w[138][160] = 5'b10000; w[138][161] = 5'b10000; w[138][162] = 5'b10000; w[138][163] = 5'b00000; w[138][164] = 5'b00000; w[138][165] = 5'b01111; w[138][166] = 5'b01111; w[138][167] = 5'b01111; w[138][168] = 5'b01111; w[138][169] = 5'b01111; w[138][170] = 5'b01111; w[138][171] = 5'b01111; w[138][172] = 5'b00000; w[138][173] = 5'b00000; w[138][174] = 5'b10000; w[138][175] = 5'b10000; w[138][176] = 5'b10000; w[138][177] = 5'b00000; w[138][178] = 5'b01111; w[138][179] = 5'b01111; w[138][180] = 5'b01111; w[138][181] = 5'b01111; w[138][182] = 5'b01111; w[138][183] = 5'b01111; w[138][184] = 5'b01111; w[138][185] = 5'b01111; w[138][186] = 5'b01111; w[138][187] = 5'b01111; w[138][188] = 5'b01111; w[138][189] = 5'b01111; w[138][190] = 5'b01111; w[138][191] = 5'b01111; w[138][192] = 5'b01111; w[138][193] = 5'b01111; w[138][194] = 5'b01111; w[138][195] = 5'b01111; w[138][196] = 5'b01111; w[138][197] = 5'b01111; w[138][198] = 5'b01111; w[138][199] = 5'b01111; w[138][200] = 5'b01111; w[138][201] = 5'b01111; w[138][202] = 5'b01111; w[138][203] = 5'b01111; w[138][204] = 5'b01111; w[138][205] = 5'b01111; w[138][206] = 5'b01111; w[138][207] = 5'b01111; w[138][208] = 5'b01111; w[138][209] = 5'b01111; 
w[139][0] = 5'b01111; w[139][1] = 5'b01111; w[139][2] = 5'b01111; w[139][3] = 5'b01111; w[139][4] = 5'b01111; w[139][5] = 5'b01111; w[139][6] = 5'b01111; w[139][7] = 5'b01111; w[139][8] = 5'b01111; w[139][9] = 5'b01111; w[139][10] = 5'b01111; w[139][11] = 5'b01111; w[139][12] = 5'b01111; w[139][13] = 5'b01111; w[139][14] = 5'b01111; w[139][15] = 5'b01111; w[139][16] = 5'b01111; w[139][17] = 5'b01111; w[139][18] = 5'b01111; w[139][19] = 5'b01111; w[139][20] = 5'b01111; w[139][21] = 5'b01111; w[139][22] = 5'b01111; w[139][23] = 5'b01111; w[139][24] = 5'b01111; w[139][25] = 5'b01111; w[139][26] = 5'b01111; w[139][27] = 5'b01111; w[139][28] = 5'b01111; w[139][29] = 5'b01111; w[139][30] = 5'b01111; w[139][31] = 5'b00000; w[139][32] = 5'b10000; w[139][33] = 5'b10000; w[139][34] = 5'b10000; w[139][35] = 5'b10000; w[139][36] = 5'b10000; w[139][37] = 5'b10000; w[139][38] = 5'b00000; w[139][39] = 5'b01111; w[139][40] = 5'b01111; w[139][41] = 5'b01111; w[139][42] = 5'b01111; w[139][43] = 5'b01111; w[139][44] = 5'b01111; w[139][45] = 5'b10000; w[139][46] = 5'b10000; w[139][47] = 5'b10000; w[139][48] = 5'b10000; w[139][49] = 5'b10000; w[139][50] = 5'b10000; w[139][51] = 5'b10000; w[139][52] = 5'b10000; w[139][53] = 5'b01111; w[139][54] = 5'b01111; w[139][55] = 5'b01111; w[139][56] = 5'b01111; w[139][57] = 5'b01111; w[139][58] = 5'b01111; w[139][59] = 5'b00000; w[139][60] = 5'b00000; w[139][61] = 5'b01111; w[139][62] = 5'b10000; w[139][63] = 5'b00000; w[139][64] = 5'b01111; w[139][65] = 5'b00000; w[139][66] = 5'b00000; w[139][67] = 5'b01111; w[139][68] = 5'b01111; w[139][69] = 5'b01111; w[139][70] = 5'b01111; w[139][71] = 5'b01111; w[139][72] = 5'b01111; w[139][73] = 5'b00000; w[139][74] = 5'b01111; w[139][75] = 5'b01111; w[139][76] = 5'b10000; w[139][77] = 5'b00000; w[139][78] = 5'b01111; w[139][79] = 5'b01111; w[139][80] = 5'b00000; w[139][81] = 5'b01111; w[139][82] = 5'b01111; w[139][83] = 5'b01111; w[139][84] = 5'b01111; w[139][85] = 5'b01111; w[139][86] = 5'b01111; w[139][87] = 5'b00000; w[139][88] = 5'b01111; w[139][89] = 5'b01111; w[139][90] = 5'b10000; w[139][91] = 5'b10000; w[139][92] = 5'b01111; w[139][93] = 5'b01111; w[139][94] = 5'b01111; w[139][95] = 5'b01111; w[139][96] = 5'b01111; w[139][97] = 5'b01111; w[139][98] = 5'b01111; w[139][99] = 5'b01111; w[139][100] = 5'b01111; w[139][101] = 5'b00000; w[139][102] = 5'b01111; w[139][103] = 5'b01111; w[139][104] = 5'b10000; w[139][105] = 5'b10000; w[139][106] = 5'b01111; w[139][107] = 5'b00000; w[139][108] = 5'b00000; w[139][109] = 5'b01111; w[139][110] = 5'b01111; w[139][111] = 5'b01111; w[139][112] = 5'b01111; w[139][113] = 5'b01111; w[139][114] = 5'b01111; w[139][115] = 5'b00000; w[139][116] = 5'b01111; w[139][117] = 5'b01111; w[139][118] = 5'b10000; w[139][119] = 5'b10000; w[139][120] = 5'b00000; w[139][121] = 5'b00000; w[139][122] = 5'b00000; w[139][123] = 5'b01111; w[139][124] = 5'b01111; w[139][125] = 5'b01111; w[139][126] = 5'b01111; w[139][127] = 5'b01111; w[139][128] = 5'b01111; w[139][129] = 5'b00000; w[139][130] = 5'b01111; w[139][131] = 5'b01111; w[139][132] = 5'b00000; w[139][133] = 5'b10000; w[139][134] = 5'b01111; w[139][135] = 5'b01111; w[139][136] = 5'b00000; w[139][137] = 5'b01111; w[139][138] = 5'b01111; w[139][139] = 5'b00000; w[139][140] = 5'b01111; w[139][141] = 5'b01111; w[139][142] = 5'b01111; w[139][143] = 5'b00000; w[139][144] = 5'b00000; w[139][145] = 5'b01111; w[139][146] = 5'b00000; w[139][147] = 5'b10000; w[139][148] = 5'b01111; w[139][149] = 5'b00000; w[139][150] = 5'b00000; w[139][151] = 5'b01111; w[139][152] = 5'b01111; w[139][153] = 5'b01111; w[139][154] = 5'b01111; w[139][155] = 5'b01111; w[139][156] = 5'b01111; w[139][157] = 5'b00000; w[139][158] = 5'b00000; w[139][159] = 5'b00000; w[139][160] = 5'b10000; w[139][161] = 5'b10000; w[139][162] = 5'b10000; w[139][163] = 5'b00000; w[139][164] = 5'b00000; w[139][165] = 5'b01111; w[139][166] = 5'b01111; w[139][167] = 5'b01111; w[139][168] = 5'b01111; w[139][169] = 5'b01111; w[139][170] = 5'b01111; w[139][171] = 5'b01111; w[139][172] = 5'b00000; w[139][173] = 5'b00000; w[139][174] = 5'b10000; w[139][175] = 5'b10000; w[139][176] = 5'b10000; w[139][177] = 5'b00000; w[139][178] = 5'b01111; w[139][179] = 5'b01111; w[139][180] = 5'b01111; w[139][181] = 5'b01111; w[139][182] = 5'b01111; w[139][183] = 5'b01111; w[139][184] = 5'b01111; w[139][185] = 5'b01111; w[139][186] = 5'b01111; w[139][187] = 5'b01111; w[139][188] = 5'b01111; w[139][189] = 5'b01111; w[139][190] = 5'b01111; w[139][191] = 5'b01111; w[139][192] = 5'b01111; w[139][193] = 5'b01111; w[139][194] = 5'b01111; w[139][195] = 5'b01111; w[139][196] = 5'b01111; w[139][197] = 5'b01111; w[139][198] = 5'b01111; w[139][199] = 5'b01111; w[139][200] = 5'b01111; w[139][201] = 5'b01111; w[139][202] = 5'b01111; w[139][203] = 5'b01111; w[139][204] = 5'b01111; w[139][205] = 5'b01111; w[139][206] = 5'b01111; w[139][207] = 5'b01111; w[139][208] = 5'b01111; w[139][209] = 5'b01111; 
w[140][0] = 5'b01111; w[140][1] = 5'b01111; w[140][2] = 5'b01111; w[140][3] = 5'b01111; w[140][4] = 5'b01111; w[140][5] = 5'b01111; w[140][6] = 5'b01111; w[140][7] = 5'b01111; w[140][8] = 5'b01111; w[140][9] = 5'b01111; w[140][10] = 5'b01111; w[140][11] = 5'b01111; w[140][12] = 5'b01111; w[140][13] = 5'b01111; w[140][14] = 5'b01111; w[140][15] = 5'b01111; w[140][16] = 5'b01111; w[140][17] = 5'b01111; w[140][18] = 5'b01111; w[140][19] = 5'b01111; w[140][20] = 5'b01111; w[140][21] = 5'b01111; w[140][22] = 5'b01111; w[140][23] = 5'b01111; w[140][24] = 5'b01111; w[140][25] = 5'b01111; w[140][26] = 5'b01111; w[140][27] = 5'b01111; w[140][28] = 5'b01111; w[140][29] = 5'b01111; w[140][30] = 5'b01111; w[140][31] = 5'b00000; w[140][32] = 5'b10000; w[140][33] = 5'b10000; w[140][34] = 5'b10000; w[140][35] = 5'b10000; w[140][36] = 5'b10000; w[140][37] = 5'b10000; w[140][38] = 5'b00000; w[140][39] = 5'b01111; w[140][40] = 5'b01111; w[140][41] = 5'b01111; w[140][42] = 5'b01111; w[140][43] = 5'b01111; w[140][44] = 5'b01111; w[140][45] = 5'b10000; w[140][46] = 5'b10000; w[140][47] = 5'b10000; w[140][48] = 5'b10000; w[140][49] = 5'b10000; w[140][50] = 5'b10000; w[140][51] = 5'b10000; w[140][52] = 5'b10000; w[140][53] = 5'b01111; w[140][54] = 5'b01111; w[140][55] = 5'b01111; w[140][56] = 5'b01111; w[140][57] = 5'b01111; w[140][58] = 5'b01111; w[140][59] = 5'b00000; w[140][60] = 5'b00000; w[140][61] = 5'b01111; w[140][62] = 5'b10000; w[140][63] = 5'b00000; w[140][64] = 5'b01111; w[140][65] = 5'b00000; w[140][66] = 5'b00000; w[140][67] = 5'b01111; w[140][68] = 5'b01111; w[140][69] = 5'b01111; w[140][70] = 5'b01111; w[140][71] = 5'b01111; w[140][72] = 5'b01111; w[140][73] = 5'b00000; w[140][74] = 5'b01111; w[140][75] = 5'b01111; w[140][76] = 5'b10000; w[140][77] = 5'b00000; w[140][78] = 5'b01111; w[140][79] = 5'b01111; w[140][80] = 5'b00000; w[140][81] = 5'b01111; w[140][82] = 5'b01111; w[140][83] = 5'b01111; w[140][84] = 5'b01111; w[140][85] = 5'b01111; w[140][86] = 5'b01111; w[140][87] = 5'b00000; w[140][88] = 5'b01111; w[140][89] = 5'b01111; w[140][90] = 5'b10000; w[140][91] = 5'b10000; w[140][92] = 5'b01111; w[140][93] = 5'b01111; w[140][94] = 5'b01111; w[140][95] = 5'b01111; w[140][96] = 5'b01111; w[140][97] = 5'b01111; w[140][98] = 5'b01111; w[140][99] = 5'b01111; w[140][100] = 5'b01111; w[140][101] = 5'b00000; w[140][102] = 5'b01111; w[140][103] = 5'b01111; w[140][104] = 5'b10000; w[140][105] = 5'b10000; w[140][106] = 5'b01111; w[140][107] = 5'b00000; w[140][108] = 5'b00000; w[140][109] = 5'b01111; w[140][110] = 5'b01111; w[140][111] = 5'b01111; w[140][112] = 5'b01111; w[140][113] = 5'b01111; w[140][114] = 5'b01111; w[140][115] = 5'b00000; w[140][116] = 5'b01111; w[140][117] = 5'b01111; w[140][118] = 5'b10000; w[140][119] = 5'b10000; w[140][120] = 5'b00000; w[140][121] = 5'b00000; w[140][122] = 5'b00000; w[140][123] = 5'b01111; w[140][124] = 5'b01111; w[140][125] = 5'b01111; w[140][126] = 5'b01111; w[140][127] = 5'b01111; w[140][128] = 5'b01111; w[140][129] = 5'b00000; w[140][130] = 5'b01111; w[140][131] = 5'b01111; w[140][132] = 5'b00000; w[140][133] = 5'b10000; w[140][134] = 5'b01111; w[140][135] = 5'b01111; w[140][136] = 5'b00000; w[140][137] = 5'b01111; w[140][138] = 5'b01111; w[140][139] = 5'b01111; w[140][140] = 5'b00000; w[140][141] = 5'b01111; w[140][142] = 5'b01111; w[140][143] = 5'b00000; w[140][144] = 5'b00000; w[140][145] = 5'b01111; w[140][146] = 5'b00000; w[140][147] = 5'b10000; w[140][148] = 5'b01111; w[140][149] = 5'b00000; w[140][150] = 5'b00000; w[140][151] = 5'b01111; w[140][152] = 5'b01111; w[140][153] = 5'b01111; w[140][154] = 5'b01111; w[140][155] = 5'b01111; w[140][156] = 5'b01111; w[140][157] = 5'b00000; w[140][158] = 5'b00000; w[140][159] = 5'b00000; w[140][160] = 5'b10000; w[140][161] = 5'b10000; w[140][162] = 5'b10000; w[140][163] = 5'b00000; w[140][164] = 5'b00000; w[140][165] = 5'b01111; w[140][166] = 5'b01111; w[140][167] = 5'b01111; w[140][168] = 5'b01111; w[140][169] = 5'b01111; w[140][170] = 5'b01111; w[140][171] = 5'b01111; w[140][172] = 5'b00000; w[140][173] = 5'b00000; w[140][174] = 5'b10000; w[140][175] = 5'b10000; w[140][176] = 5'b10000; w[140][177] = 5'b00000; w[140][178] = 5'b01111; w[140][179] = 5'b01111; w[140][180] = 5'b01111; w[140][181] = 5'b01111; w[140][182] = 5'b01111; w[140][183] = 5'b01111; w[140][184] = 5'b01111; w[140][185] = 5'b01111; w[140][186] = 5'b01111; w[140][187] = 5'b01111; w[140][188] = 5'b01111; w[140][189] = 5'b01111; w[140][190] = 5'b01111; w[140][191] = 5'b01111; w[140][192] = 5'b01111; w[140][193] = 5'b01111; w[140][194] = 5'b01111; w[140][195] = 5'b01111; w[140][196] = 5'b01111; w[140][197] = 5'b01111; w[140][198] = 5'b01111; w[140][199] = 5'b01111; w[140][200] = 5'b01111; w[140][201] = 5'b01111; w[140][202] = 5'b01111; w[140][203] = 5'b01111; w[140][204] = 5'b01111; w[140][205] = 5'b01111; w[140][206] = 5'b01111; w[140][207] = 5'b01111; w[140][208] = 5'b01111; w[140][209] = 5'b01111; 
w[141][0] = 5'b01111; w[141][1] = 5'b01111; w[141][2] = 5'b01111; w[141][3] = 5'b01111; w[141][4] = 5'b01111; w[141][5] = 5'b01111; w[141][6] = 5'b01111; w[141][7] = 5'b01111; w[141][8] = 5'b01111; w[141][9] = 5'b01111; w[141][10] = 5'b01111; w[141][11] = 5'b01111; w[141][12] = 5'b01111; w[141][13] = 5'b01111; w[141][14] = 5'b01111; w[141][15] = 5'b01111; w[141][16] = 5'b01111; w[141][17] = 5'b01111; w[141][18] = 5'b01111; w[141][19] = 5'b01111; w[141][20] = 5'b01111; w[141][21] = 5'b01111; w[141][22] = 5'b01111; w[141][23] = 5'b01111; w[141][24] = 5'b01111; w[141][25] = 5'b01111; w[141][26] = 5'b01111; w[141][27] = 5'b01111; w[141][28] = 5'b01111; w[141][29] = 5'b01111; w[141][30] = 5'b01111; w[141][31] = 5'b00000; w[141][32] = 5'b10000; w[141][33] = 5'b10000; w[141][34] = 5'b10000; w[141][35] = 5'b10000; w[141][36] = 5'b10000; w[141][37] = 5'b10000; w[141][38] = 5'b00000; w[141][39] = 5'b01111; w[141][40] = 5'b01111; w[141][41] = 5'b01111; w[141][42] = 5'b01111; w[141][43] = 5'b01111; w[141][44] = 5'b01111; w[141][45] = 5'b10000; w[141][46] = 5'b10000; w[141][47] = 5'b10000; w[141][48] = 5'b10000; w[141][49] = 5'b10000; w[141][50] = 5'b10000; w[141][51] = 5'b10000; w[141][52] = 5'b10000; w[141][53] = 5'b01111; w[141][54] = 5'b01111; w[141][55] = 5'b01111; w[141][56] = 5'b01111; w[141][57] = 5'b01111; w[141][58] = 5'b01111; w[141][59] = 5'b00000; w[141][60] = 5'b00000; w[141][61] = 5'b01111; w[141][62] = 5'b10000; w[141][63] = 5'b00000; w[141][64] = 5'b01111; w[141][65] = 5'b00000; w[141][66] = 5'b00000; w[141][67] = 5'b01111; w[141][68] = 5'b01111; w[141][69] = 5'b01111; w[141][70] = 5'b01111; w[141][71] = 5'b01111; w[141][72] = 5'b01111; w[141][73] = 5'b00000; w[141][74] = 5'b01111; w[141][75] = 5'b01111; w[141][76] = 5'b10000; w[141][77] = 5'b00000; w[141][78] = 5'b01111; w[141][79] = 5'b01111; w[141][80] = 5'b00000; w[141][81] = 5'b01111; w[141][82] = 5'b01111; w[141][83] = 5'b01111; w[141][84] = 5'b01111; w[141][85] = 5'b01111; w[141][86] = 5'b01111; w[141][87] = 5'b00000; w[141][88] = 5'b01111; w[141][89] = 5'b01111; w[141][90] = 5'b10000; w[141][91] = 5'b10000; w[141][92] = 5'b01111; w[141][93] = 5'b01111; w[141][94] = 5'b01111; w[141][95] = 5'b01111; w[141][96] = 5'b01111; w[141][97] = 5'b01111; w[141][98] = 5'b01111; w[141][99] = 5'b01111; w[141][100] = 5'b01111; w[141][101] = 5'b00000; w[141][102] = 5'b01111; w[141][103] = 5'b01111; w[141][104] = 5'b10000; w[141][105] = 5'b10000; w[141][106] = 5'b01111; w[141][107] = 5'b00000; w[141][108] = 5'b00000; w[141][109] = 5'b01111; w[141][110] = 5'b01111; w[141][111] = 5'b01111; w[141][112] = 5'b01111; w[141][113] = 5'b01111; w[141][114] = 5'b01111; w[141][115] = 5'b00000; w[141][116] = 5'b01111; w[141][117] = 5'b01111; w[141][118] = 5'b10000; w[141][119] = 5'b10000; w[141][120] = 5'b00000; w[141][121] = 5'b00000; w[141][122] = 5'b00000; w[141][123] = 5'b01111; w[141][124] = 5'b01111; w[141][125] = 5'b01111; w[141][126] = 5'b01111; w[141][127] = 5'b01111; w[141][128] = 5'b01111; w[141][129] = 5'b00000; w[141][130] = 5'b01111; w[141][131] = 5'b01111; w[141][132] = 5'b00000; w[141][133] = 5'b10000; w[141][134] = 5'b01111; w[141][135] = 5'b01111; w[141][136] = 5'b00000; w[141][137] = 5'b01111; w[141][138] = 5'b01111; w[141][139] = 5'b01111; w[141][140] = 5'b01111; w[141][141] = 5'b00000; w[141][142] = 5'b01111; w[141][143] = 5'b00000; w[141][144] = 5'b00000; w[141][145] = 5'b01111; w[141][146] = 5'b00000; w[141][147] = 5'b10000; w[141][148] = 5'b01111; w[141][149] = 5'b00000; w[141][150] = 5'b00000; w[141][151] = 5'b01111; w[141][152] = 5'b01111; w[141][153] = 5'b01111; w[141][154] = 5'b01111; w[141][155] = 5'b01111; w[141][156] = 5'b01111; w[141][157] = 5'b00000; w[141][158] = 5'b00000; w[141][159] = 5'b00000; w[141][160] = 5'b10000; w[141][161] = 5'b10000; w[141][162] = 5'b10000; w[141][163] = 5'b00000; w[141][164] = 5'b00000; w[141][165] = 5'b01111; w[141][166] = 5'b01111; w[141][167] = 5'b01111; w[141][168] = 5'b01111; w[141][169] = 5'b01111; w[141][170] = 5'b01111; w[141][171] = 5'b01111; w[141][172] = 5'b00000; w[141][173] = 5'b00000; w[141][174] = 5'b10000; w[141][175] = 5'b10000; w[141][176] = 5'b10000; w[141][177] = 5'b00000; w[141][178] = 5'b01111; w[141][179] = 5'b01111; w[141][180] = 5'b01111; w[141][181] = 5'b01111; w[141][182] = 5'b01111; w[141][183] = 5'b01111; w[141][184] = 5'b01111; w[141][185] = 5'b01111; w[141][186] = 5'b01111; w[141][187] = 5'b01111; w[141][188] = 5'b01111; w[141][189] = 5'b01111; w[141][190] = 5'b01111; w[141][191] = 5'b01111; w[141][192] = 5'b01111; w[141][193] = 5'b01111; w[141][194] = 5'b01111; w[141][195] = 5'b01111; w[141][196] = 5'b01111; w[141][197] = 5'b01111; w[141][198] = 5'b01111; w[141][199] = 5'b01111; w[141][200] = 5'b01111; w[141][201] = 5'b01111; w[141][202] = 5'b01111; w[141][203] = 5'b01111; w[141][204] = 5'b01111; w[141][205] = 5'b01111; w[141][206] = 5'b01111; w[141][207] = 5'b01111; w[141][208] = 5'b01111; w[141][209] = 5'b01111; 
w[142][0] = 5'b01111; w[142][1] = 5'b01111; w[142][2] = 5'b01111; w[142][3] = 5'b01111; w[142][4] = 5'b01111; w[142][5] = 5'b01111; w[142][6] = 5'b01111; w[142][7] = 5'b01111; w[142][8] = 5'b01111; w[142][9] = 5'b01111; w[142][10] = 5'b01111; w[142][11] = 5'b01111; w[142][12] = 5'b01111; w[142][13] = 5'b01111; w[142][14] = 5'b01111; w[142][15] = 5'b01111; w[142][16] = 5'b01111; w[142][17] = 5'b01111; w[142][18] = 5'b01111; w[142][19] = 5'b01111; w[142][20] = 5'b01111; w[142][21] = 5'b01111; w[142][22] = 5'b01111; w[142][23] = 5'b01111; w[142][24] = 5'b01111; w[142][25] = 5'b01111; w[142][26] = 5'b01111; w[142][27] = 5'b01111; w[142][28] = 5'b01111; w[142][29] = 5'b01111; w[142][30] = 5'b00000; w[142][31] = 5'b10000; w[142][32] = 5'b00000; w[142][33] = 5'b10000; w[142][34] = 5'b00000; w[142][35] = 5'b00000; w[142][36] = 5'b00000; w[142][37] = 5'b00000; w[142][38] = 5'b10000; w[142][39] = 5'b00000; w[142][40] = 5'b01111; w[142][41] = 5'b01111; w[142][42] = 5'b01111; w[142][43] = 5'b01111; w[142][44] = 5'b00000; w[142][45] = 5'b00000; w[142][46] = 5'b00000; w[142][47] = 5'b10000; w[142][48] = 5'b00000; w[142][49] = 5'b00000; w[142][50] = 5'b00000; w[142][51] = 5'b00000; w[142][52] = 5'b00000; w[142][53] = 5'b00000; w[142][54] = 5'b01111; w[142][55] = 5'b01111; w[142][56] = 5'b01111; w[142][57] = 5'b01111; w[142][58] = 5'b01111; w[142][59] = 5'b01111; w[142][60] = 5'b01111; w[142][61] = 5'b00000; w[142][62] = 5'b10000; w[142][63] = 5'b10000; w[142][64] = 5'b01111; w[142][65] = 5'b01111; w[142][66] = 5'b01111; w[142][67] = 5'b01111; w[142][68] = 5'b01111; w[142][69] = 5'b01111; w[142][70] = 5'b01111; w[142][71] = 5'b01111; w[142][72] = 5'b01111; w[142][73] = 5'b01111; w[142][74] = 5'b00000; w[142][75] = 5'b00000; w[142][76] = 5'b10000; w[142][77] = 5'b10000; w[142][78] = 5'b01111; w[142][79] = 5'b00000; w[142][80] = 5'b01111; w[142][81] = 5'b01111; w[142][82] = 5'b01111; w[142][83] = 5'b01111; w[142][84] = 5'b01111; w[142][85] = 5'b01111; w[142][86] = 5'b01111; w[142][87] = 5'b01111; w[142][88] = 5'b00000; w[142][89] = 5'b00000; w[142][90] = 5'b10000; w[142][91] = 5'b10000; w[142][92] = 5'b01111; w[142][93] = 5'b00000; w[142][94] = 5'b00000; w[142][95] = 5'b01111; w[142][96] = 5'b01111; w[142][97] = 5'b01111; w[142][98] = 5'b01111; w[142][99] = 5'b01111; w[142][100] = 5'b01111; w[142][101] = 5'b01111; w[142][102] = 5'b00000; w[142][103] = 5'b01111; w[142][104] = 5'b10000; w[142][105] = 5'b10000; w[142][106] = 5'b01111; w[142][107] = 5'b01111; w[142][108] = 5'b01111; w[142][109] = 5'b01111; w[142][110] = 5'b01111; w[142][111] = 5'b01111; w[142][112] = 5'b01111; w[142][113] = 5'b01111; w[142][114] = 5'b01111; w[142][115] = 5'b01111; w[142][116] = 5'b00000; w[142][117] = 5'b01111; w[142][118] = 5'b10000; w[142][119] = 5'b10000; w[142][120] = 5'b01111; w[142][121] = 5'b01111; w[142][122] = 5'b01111; w[142][123] = 5'b01111; w[142][124] = 5'b01111; w[142][125] = 5'b01111; w[142][126] = 5'b01111; w[142][127] = 5'b01111; w[142][128] = 5'b01111; w[142][129] = 5'b01111; w[142][130] = 5'b00000; w[142][131] = 5'b01111; w[142][132] = 5'b10000; w[142][133] = 5'b10000; w[142][134] = 5'b00000; w[142][135] = 5'b00000; w[142][136] = 5'b01111; w[142][137] = 5'b01111; w[142][138] = 5'b01111; w[142][139] = 5'b01111; w[142][140] = 5'b01111; w[142][141] = 5'b01111; w[142][142] = 5'b00000; w[142][143] = 5'b01111; w[142][144] = 5'b01111; w[142][145] = 5'b01111; w[142][146] = 5'b10000; w[142][147] = 5'b10000; w[142][148] = 5'b00000; w[142][149] = 5'b01111; w[142][150] = 5'b01111; w[142][151] = 5'b01111; w[142][152] = 5'b01111; w[142][153] = 5'b01111; w[142][154] = 5'b01111; w[142][155] = 5'b01111; w[142][156] = 5'b01111; w[142][157] = 5'b01111; w[142][158] = 5'b01111; w[142][159] = 5'b01111; w[142][160] = 5'b00000; w[142][161] = 5'b00000; w[142][162] = 5'b00000; w[142][163] = 5'b01111; w[142][164] = 5'b01111; w[142][165] = 5'b01111; w[142][166] = 5'b01111; w[142][167] = 5'b01111; w[142][168] = 5'b01111; w[142][169] = 5'b01111; w[142][170] = 5'b01111; w[142][171] = 5'b00000; w[142][172] = 5'b01111; w[142][173] = 5'b01111; w[142][174] = 5'b00000; w[142][175] = 5'b00000; w[142][176] = 5'b00000; w[142][177] = 5'b01111; w[142][178] = 5'b00000; w[142][179] = 5'b01111; w[142][180] = 5'b01111; w[142][181] = 5'b01111; w[142][182] = 5'b01111; w[142][183] = 5'b01111; w[142][184] = 5'b01111; w[142][185] = 5'b01111; w[142][186] = 5'b01111; w[142][187] = 5'b01111; w[142][188] = 5'b01111; w[142][189] = 5'b01111; w[142][190] = 5'b01111; w[142][191] = 5'b01111; w[142][192] = 5'b01111; w[142][193] = 5'b01111; w[142][194] = 5'b01111; w[142][195] = 5'b01111; w[142][196] = 5'b01111; w[142][197] = 5'b01111; w[142][198] = 5'b01111; w[142][199] = 5'b01111; w[142][200] = 5'b01111; w[142][201] = 5'b01111; w[142][202] = 5'b01111; w[142][203] = 5'b01111; w[142][204] = 5'b01111; w[142][205] = 5'b01111; w[142][206] = 5'b01111; w[142][207] = 5'b01111; w[142][208] = 5'b01111; w[142][209] = 5'b01111; 
w[143][0] = 5'b00000; w[143][1] = 5'b00000; w[143][2] = 5'b00000; w[143][3] = 5'b00000; w[143][4] = 5'b00000; w[143][5] = 5'b00000; w[143][6] = 5'b00000; w[143][7] = 5'b00000; w[143][8] = 5'b00000; w[143][9] = 5'b00000; w[143][10] = 5'b00000; w[143][11] = 5'b00000; w[143][12] = 5'b00000; w[143][13] = 5'b00000; w[143][14] = 5'b00000; w[143][15] = 5'b00000; w[143][16] = 5'b00000; w[143][17] = 5'b00000; w[143][18] = 5'b00000; w[143][19] = 5'b00000; w[143][20] = 5'b00000; w[143][21] = 5'b00000; w[143][22] = 5'b00000; w[143][23] = 5'b00000; w[143][24] = 5'b00000; w[143][25] = 5'b00000; w[143][26] = 5'b00000; w[143][27] = 5'b00000; w[143][28] = 5'b00000; w[143][29] = 5'b00000; w[143][30] = 5'b10000; w[143][31] = 5'b00000; w[143][32] = 5'b01111; w[143][33] = 5'b00000; w[143][34] = 5'b10000; w[143][35] = 5'b10000; w[143][36] = 5'b10000; w[143][37] = 5'b01111; w[143][38] = 5'b00000; w[143][39] = 5'b10000; w[143][40] = 5'b00000; w[143][41] = 5'b00000; w[143][42] = 5'b00000; w[143][43] = 5'b00000; w[143][44] = 5'b10000; w[143][45] = 5'b01111; w[143][46] = 5'b01111; w[143][47] = 5'b00000; w[143][48] = 5'b10000; w[143][49] = 5'b10000; w[143][50] = 5'b10000; w[143][51] = 5'b01111; w[143][52] = 5'b01111; w[143][53] = 5'b10000; w[143][54] = 5'b00000; w[143][55] = 5'b00000; w[143][56] = 5'b00000; w[143][57] = 5'b00000; w[143][58] = 5'b01111; w[143][59] = 5'b01111; w[143][60] = 5'b01111; w[143][61] = 5'b01111; w[143][62] = 5'b10000; w[143][63] = 5'b10000; w[143][64] = 5'b00000; w[143][65] = 5'b01111; w[143][66] = 5'b01111; w[143][67] = 5'b01111; w[143][68] = 5'b00000; w[143][69] = 5'b00000; w[143][70] = 5'b00000; w[143][71] = 5'b00000; w[143][72] = 5'b01111; w[143][73] = 5'b01111; w[143][74] = 5'b01111; w[143][75] = 5'b01111; w[143][76] = 5'b10000; w[143][77] = 5'b10000; w[143][78] = 5'b00000; w[143][79] = 5'b01111; w[143][80] = 5'b01111; w[143][81] = 5'b01111; w[143][82] = 5'b00000; w[143][83] = 5'b00000; w[143][84] = 5'b00000; w[143][85] = 5'b00000; w[143][86] = 5'b01111; w[143][87] = 5'b01111; w[143][88] = 5'b01111; w[143][89] = 5'b01111; w[143][90] = 5'b10000; w[143][91] = 5'b10000; w[143][92] = 5'b00000; w[143][93] = 5'b01111; w[143][94] = 5'b01111; w[143][95] = 5'b00000; w[143][96] = 5'b00000; w[143][97] = 5'b00000; w[143][98] = 5'b00000; w[143][99] = 5'b00000; w[143][100] = 5'b01111; w[143][101] = 5'b01111; w[143][102] = 5'b01111; w[143][103] = 5'b00000; w[143][104] = 5'b10000; w[143][105] = 5'b10000; w[143][106] = 5'b01111; w[143][107] = 5'b01111; w[143][108] = 5'b01111; w[143][109] = 5'b01111; w[143][110] = 5'b00000; w[143][111] = 5'b00000; w[143][112] = 5'b00000; w[143][113] = 5'b00000; w[143][114] = 5'b01111; w[143][115] = 5'b01111; w[143][116] = 5'b01111; w[143][117] = 5'b00000; w[143][118] = 5'b10000; w[143][119] = 5'b10000; w[143][120] = 5'b01111; w[143][121] = 5'b01111; w[143][122] = 5'b01111; w[143][123] = 5'b01111; w[143][124] = 5'b00000; w[143][125] = 5'b00000; w[143][126] = 5'b00000; w[143][127] = 5'b00000; w[143][128] = 5'b01111; w[143][129] = 5'b01111; w[143][130] = 5'b01111; w[143][131] = 5'b00000; w[143][132] = 5'b10000; w[143][133] = 5'b10000; w[143][134] = 5'b01111; w[143][135] = 5'b01111; w[143][136] = 5'b01111; w[143][137] = 5'b01111; w[143][138] = 5'b00000; w[143][139] = 5'b00000; w[143][140] = 5'b00000; w[143][141] = 5'b00000; w[143][142] = 5'b01111; w[143][143] = 5'b00000; w[143][144] = 5'b01111; w[143][145] = 5'b00000; w[143][146] = 5'b10000; w[143][147] = 5'b10000; w[143][148] = 5'b01111; w[143][149] = 5'b01111; w[143][150] = 5'b01111; w[143][151] = 5'b01111; w[143][152] = 5'b00000; w[143][153] = 5'b00000; w[143][154] = 5'b00000; w[143][155] = 5'b00000; w[143][156] = 5'b00000; w[143][157] = 5'b01111; w[143][158] = 5'b01111; w[143][159] = 5'b00000; w[143][160] = 5'b10000; w[143][161] = 5'b10000; w[143][162] = 5'b01111; w[143][163] = 5'b01111; w[143][164] = 5'b01111; w[143][165] = 5'b00000; w[143][166] = 5'b00000; w[143][167] = 5'b00000; w[143][168] = 5'b00000; w[143][169] = 5'b00000; w[143][170] = 5'b00000; w[143][171] = 5'b01111; w[143][172] = 5'b01111; w[143][173] = 5'b00000; w[143][174] = 5'b10000; w[143][175] = 5'b10000; w[143][176] = 5'b01111; w[143][177] = 5'b01111; w[143][178] = 5'b01111; w[143][179] = 5'b00000; w[143][180] = 5'b00000; w[143][181] = 5'b00000; w[143][182] = 5'b00000; w[143][183] = 5'b00000; w[143][184] = 5'b00000; w[143][185] = 5'b00000; w[143][186] = 5'b00000; w[143][187] = 5'b00000; w[143][188] = 5'b00000; w[143][189] = 5'b00000; w[143][190] = 5'b00000; w[143][191] = 5'b00000; w[143][192] = 5'b00000; w[143][193] = 5'b00000; w[143][194] = 5'b00000; w[143][195] = 5'b00000; w[143][196] = 5'b00000; w[143][197] = 5'b00000; w[143][198] = 5'b00000; w[143][199] = 5'b00000; w[143][200] = 5'b00000; w[143][201] = 5'b00000; w[143][202] = 5'b00000; w[143][203] = 5'b00000; w[143][204] = 5'b00000; w[143][205] = 5'b00000; w[143][206] = 5'b00000; w[143][207] = 5'b00000; w[143][208] = 5'b00000; w[143][209] = 5'b00000; 
w[144][0] = 5'b00000; w[144][1] = 5'b00000; w[144][2] = 5'b00000; w[144][3] = 5'b00000; w[144][4] = 5'b00000; w[144][5] = 5'b00000; w[144][6] = 5'b00000; w[144][7] = 5'b00000; w[144][8] = 5'b00000; w[144][9] = 5'b00000; w[144][10] = 5'b00000; w[144][11] = 5'b00000; w[144][12] = 5'b00000; w[144][13] = 5'b00000; w[144][14] = 5'b00000; w[144][15] = 5'b00000; w[144][16] = 5'b00000; w[144][17] = 5'b00000; w[144][18] = 5'b00000; w[144][19] = 5'b00000; w[144][20] = 5'b00000; w[144][21] = 5'b00000; w[144][22] = 5'b00000; w[144][23] = 5'b00000; w[144][24] = 5'b00000; w[144][25] = 5'b00000; w[144][26] = 5'b00000; w[144][27] = 5'b00000; w[144][28] = 5'b00000; w[144][29] = 5'b00000; w[144][30] = 5'b10000; w[144][31] = 5'b00000; w[144][32] = 5'b01111; w[144][33] = 5'b00000; w[144][34] = 5'b10000; w[144][35] = 5'b10000; w[144][36] = 5'b10000; w[144][37] = 5'b01111; w[144][38] = 5'b00000; w[144][39] = 5'b10000; w[144][40] = 5'b00000; w[144][41] = 5'b00000; w[144][42] = 5'b00000; w[144][43] = 5'b00000; w[144][44] = 5'b10000; w[144][45] = 5'b01111; w[144][46] = 5'b01111; w[144][47] = 5'b00000; w[144][48] = 5'b10000; w[144][49] = 5'b10000; w[144][50] = 5'b10000; w[144][51] = 5'b01111; w[144][52] = 5'b01111; w[144][53] = 5'b10000; w[144][54] = 5'b00000; w[144][55] = 5'b00000; w[144][56] = 5'b00000; w[144][57] = 5'b00000; w[144][58] = 5'b01111; w[144][59] = 5'b01111; w[144][60] = 5'b01111; w[144][61] = 5'b01111; w[144][62] = 5'b10000; w[144][63] = 5'b10000; w[144][64] = 5'b00000; w[144][65] = 5'b01111; w[144][66] = 5'b01111; w[144][67] = 5'b01111; w[144][68] = 5'b00000; w[144][69] = 5'b00000; w[144][70] = 5'b00000; w[144][71] = 5'b00000; w[144][72] = 5'b01111; w[144][73] = 5'b01111; w[144][74] = 5'b01111; w[144][75] = 5'b01111; w[144][76] = 5'b10000; w[144][77] = 5'b10000; w[144][78] = 5'b00000; w[144][79] = 5'b01111; w[144][80] = 5'b01111; w[144][81] = 5'b01111; w[144][82] = 5'b00000; w[144][83] = 5'b00000; w[144][84] = 5'b00000; w[144][85] = 5'b00000; w[144][86] = 5'b01111; w[144][87] = 5'b01111; w[144][88] = 5'b01111; w[144][89] = 5'b01111; w[144][90] = 5'b10000; w[144][91] = 5'b10000; w[144][92] = 5'b00000; w[144][93] = 5'b01111; w[144][94] = 5'b01111; w[144][95] = 5'b00000; w[144][96] = 5'b00000; w[144][97] = 5'b00000; w[144][98] = 5'b00000; w[144][99] = 5'b00000; w[144][100] = 5'b01111; w[144][101] = 5'b01111; w[144][102] = 5'b01111; w[144][103] = 5'b00000; w[144][104] = 5'b10000; w[144][105] = 5'b10000; w[144][106] = 5'b01111; w[144][107] = 5'b01111; w[144][108] = 5'b01111; w[144][109] = 5'b01111; w[144][110] = 5'b00000; w[144][111] = 5'b00000; w[144][112] = 5'b00000; w[144][113] = 5'b00000; w[144][114] = 5'b01111; w[144][115] = 5'b01111; w[144][116] = 5'b01111; w[144][117] = 5'b00000; w[144][118] = 5'b10000; w[144][119] = 5'b10000; w[144][120] = 5'b01111; w[144][121] = 5'b01111; w[144][122] = 5'b01111; w[144][123] = 5'b01111; w[144][124] = 5'b00000; w[144][125] = 5'b00000; w[144][126] = 5'b00000; w[144][127] = 5'b00000; w[144][128] = 5'b01111; w[144][129] = 5'b01111; w[144][130] = 5'b01111; w[144][131] = 5'b00000; w[144][132] = 5'b10000; w[144][133] = 5'b10000; w[144][134] = 5'b01111; w[144][135] = 5'b01111; w[144][136] = 5'b01111; w[144][137] = 5'b01111; w[144][138] = 5'b00000; w[144][139] = 5'b00000; w[144][140] = 5'b00000; w[144][141] = 5'b00000; w[144][142] = 5'b01111; w[144][143] = 5'b01111; w[144][144] = 5'b00000; w[144][145] = 5'b00000; w[144][146] = 5'b10000; w[144][147] = 5'b10000; w[144][148] = 5'b01111; w[144][149] = 5'b01111; w[144][150] = 5'b01111; w[144][151] = 5'b01111; w[144][152] = 5'b00000; w[144][153] = 5'b00000; w[144][154] = 5'b00000; w[144][155] = 5'b00000; w[144][156] = 5'b00000; w[144][157] = 5'b01111; w[144][158] = 5'b01111; w[144][159] = 5'b00000; w[144][160] = 5'b10000; w[144][161] = 5'b10000; w[144][162] = 5'b01111; w[144][163] = 5'b01111; w[144][164] = 5'b01111; w[144][165] = 5'b00000; w[144][166] = 5'b00000; w[144][167] = 5'b00000; w[144][168] = 5'b00000; w[144][169] = 5'b00000; w[144][170] = 5'b00000; w[144][171] = 5'b01111; w[144][172] = 5'b01111; w[144][173] = 5'b00000; w[144][174] = 5'b10000; w[144][175] = 5'b10000; w[144][176] = 5'b01111; w[144][177] = 5'b01111; w[144][178] = 5'b01111; w[144][179] = 5'b00000; w[144][180] = 5'b00000; w[144][181] = 5'b00000; w[144][182] = 5'b00000; w[144][183] = 5'b00000; w[144][184] = 5'b00000; w[144][185] = 5'b00000; w[144][186] = 5'b00000; w[144][187] = 5'b00000; w[144][188] = 5'b00000; w[144][189] = 5'b00000; w[144][190] = 5'b00000; w[144][191] = 5'b00000; w[144][192] = 5'b00000; w[144][193] = 5'b00000; w[144][194] = 5'b00000; w[144][195] = 5'b00000; w[144][196] = 5'b00000; w[144][197] = 5'b00000; w[144][198] = 5'b00000; w[144][199] = 5'b00000; w[144][200] = 5'b00000; w[144][201] = 5'b00000; w[144][202] = 5'b00000; w[144][203] = 5'b00000; w[144][204] = 5'b00000; w[144][205] = 5'b00000; w[144][206] = 5'b00000; w[144][207] = 5'b00000; w[144][208] = 5'b00000; w[144][209] = 5'b00000; 
w[145][0] = 5'b01111; w[145][1] = 5'b01111; w[145][2] = 5'b01111; w[145][3] = 5'b01111; w[145][4] = 5'b01111; w[145][5] = 5'b01111; w[145][6] = 5'b01111; w[145][7] = 5'b01111; w[145][8] = 5'b01111; w[145][9] = 5'b01111; w[145][10] = 5'b01111; w[145][11] = 5'b01111; w[145][12] = 5'b01111; w[145][13] = 5'b01111; w[145][14] = 5'b01111; w[145][15] = 5'b01111; w[145][16] = 5'b01111; w[145][17] = 5'b01111; w[145][18] = 5'b01111; w[145][19] = 5'b01111; w[145][20] = 5'b01111; w[145][21] = 5'b01111; w[145][22] = 5'b01111; w[145][23] = 5'b01111; w[145][24] = 5'b01111; w[145][25] = 5'b01111; w[145][26] = 5'b01111; w[145][27] = 5'b01111; w[145][28] = 5'b01111; w[145][29] = 5'b01111; w[145][30] = 5'b01111; w[145][31] = 5'b00000; w[145][32] = 5'b10000; w[145][33] = 5'b10000; w[145][34] = 5'b10000; w[145][35] = 5'b10000; w[145][36] = 5'b10000; w[145][37] = 5'b10000; w[145][38] = 5'b00000; w[145][39] = 5'b01111; w[145][40] = 5'b01111; w[145][41] = 5'b01111; w[145][42] = 5'b01111; w[145][43] = 5'b01111; w[145][44] = 5'b01111; w[145][45] = 5'b10000; w[145][46] = 5'b10000; w[145][47] = 5'b10000; w[145][48] = 5'b10000; w[145][49] = 5'b10000; w[145][50] = 5'b10000; w[145][51] = 5'b10000; w[145][52] = 5'b10000; w[145][53] = 5'b01111; w[145][54] = 5'b01111; w[145][55] = 5'b01111; w[145][56] = 5'b01111; w[145][57] = 5'b01111; w[145][58] = 5'b01111; w[145][59] = 5'b00000; w[145][60] = 5'b00000; w[145][61] = 5'b01111; w[145][62] = 5'b10000; w[145][63] = 5'b00000; w[145][64] = 5'b01111; w[145][65] = 5'b00000; w[145][66] = 5'b00000; w[145][67] = 5'b01111; w[145][68] = 5'b01111; w[145][69] = 5'b01111; w[145][70] = 5'b01111; w[145][71] = 5'b01111; w[145][72] = 5'b01111; w[145][73] = 5'b00000; w[145][74] = 5'b01111; w[145][75] = 5'b01111; w[145][76] = 5'b10000; w[145][77] = 5'b00000; w[145][78] = 5'b01111; w[145][79] = 5'b01111; w[145][80] = 5'b00000; w[145][81] = 5'b01111; w[145][82] = 5'b01111; w[145][83] = 5'b01111; w[145][84] = 5'b01111; w[145][85] = 5'b01111; w[145][86] = 5'b01111; w[145][87] = 5'b00000; w[145][88] = 5'b01111; w[145][89] = 5'b01111; w[145][90] = 5'b10000; w[145][91] = 5'b10000; w[145][92] = 5'b01111; w[145][93] = 5'b01111; w[145][94] = 5'b01111; w[145][95] = 5'b01111; w[145][96] = 5'b01111; w[145][97] = 5'b01111; w[145][98] = 5'b01111; w[145][99] = 5'b01111; w[145][100] = 5'b01111; w[145][101] = 5'b00000; w[145][102] = 5'b01111; w[145][103] = 5'b01111; w[145][104] = 5'b10000; w[145][105] = 5'b10000; w[145][106] = 5'b01111; w[145][107] = 5'b00000; w[145][108] = 5'b00000; w[145][109] = 5'b01111; w[145][110] = 5'b01111; w[145][111] = 5'b01111; w[145][112] = 5'b01111; w[145][113] = 5'b01111; w[145][114] = 5'b01111; w[145][115] = 5'b00000; w[145][116] = 5'b01111; w[145][117] = 5'b01111; w[145][118] = 5'b10000; w[145][119] = 5'b10000; w[145][120] = 5'b00000; w[145][121] = 5'b00000; w[145][122] = 5'b00000; w[145][123] = 5'b01111; w[145][124] = 5'b01111; w[145][125] = 5'b01111; w[145][126] = 5'b01111; w[145][127] = 5'b01111; w[145][128] = 5'b01111; w[145][129] = 5'b00000; w[145][130] = 5'b01111; w[145][131] = 5'b01111; w[145][132] = 5'b00000; w[145][133] = 5'b10000; w[145][134] = 5'b01111; w[145][135] = 5'b01111; w[145][136] = 5'b00000; w[145][137] = 5'b01111; w[145][138] = 5'b01111; w[145][139] = 5'b01111; w[145][140] = 5'b01111; w[145][141] = 5'b01111; w[145][142] = 5'b01111; w[145][143] = 5'b00000; w[145][144] = 5'b00000; w[145][145] = 5'b00000; w[145][146] = 5'b00000; w[145][147] = 5'b10000; w[145][148] = 5'b01111; w[145][149] = 5'b00000; w[145][150] = 5'b00000; w[145][151] = 5'b01111; w[145][152] = 5'b01111; w[145][153] = 5'b01111; w[145][154] = 5'b01111; w[145][155] = 5'b01111; w[145][156] = 5'b01111; w[145][157] = 5'b00000; w[145][158] = 5'b00000; w[145][159] = 5'b00000; w[145][160] = 5'b10000; w[145][161] = 5'b10000; w[145][162] = 5'b10000; w[145][163] = 5'b00000; w[145][164] = 5'b00000; w[145][165] = 5'b01111; w[145][166] = 5'b01111; w[145][167] = 5'b01111; w[145][168] = 5'b01111; w[145][169] = 5'b01111; w[145][170] = 5'b01111; w[145][171] = 5'b01111; w[145][172] = 5'b00000; w[145][173] = 5'b00000; w[145][174] = 5'b10000; w[145][175] = 5'b10000; w[145][176] = 5'b10000; w[145][177] = 5'b00000; w[145][178] = 5'b01111; w[145][179] = 5'b01111; w[145][180] = 5'b01111; w[145][181] = 5'b01111; w[145][182] = 5'b01111; w[145][183] = 5'b01111; w[145][184] = 5'b01111; w[145][185] = 5'b01111; w[145][186] = 5'b01111; w[145][187] = 5'b01111; w[145][188] = 5'b01111; w[145][189] = 5'b01111; w[145][190] = 5'b01111; w[145][191] = 5'b01111; w[145][192] = 5'b01111; w[145][193] = 5'b01111; w[145][194] = 5'b01111; w[145][195] = 5'b01111; w[145][196] = 5'b01111; w[145][197] = 5'b01111; w[145][198] = 5'b01111; w[145][199] = 5'b01111; w[145][200] = 5'b01111; w[145][201] = 5'b01111; w[145][202] = 5'b01111; w[145][203] = 5'b01111; w[145][204] = 5'b01111; w[145][205] = 5'b01111; w[145][206] = 5'b01111; w[145][207] = 5'b01111; w[145][208] = 5'b01111; w[145][209] = 5'b01111; 
w[146][0] = 5'b00000; w[146][1] = 5'b00000; w[146][2] = 5'b00000; w[146][3] = 5'b00000; w[146][4] = 5'b00000; w[146][5] = 5'b00000; w[146][6] = 5'b00000; w[146][7] = 5'b00000; w[146][8] = 5'b00000; w[146][9] = 5'b00000; w[146][10] = 5'b00000; w[146][11] = 5'b00000; w[146][12] = 5'b00000; w[146][13] = 5'b00000; w[146][14] = 5'b00000; w[146][15] = 5'b00000; w[146][16] = 5'b00000; w[146][17] = 5'b00000; w[146][18] = 5'b00000; w[146][19] = 5'b00000; w[146][20] = 5'b00000; w[146][21] = 5'b00000; w[146][22] = 5'b00000; w[146][23] = 5'b00000; w[146][24] = 5'b00000; w[146][25] = 5'b00000; w[146][26] = 5'b00000; w[146][27] = 5'b00000; w[146][28] = 5'b00000; w[146][29] = 5'b00000; w[146][30] = 5'b01111; w[146][31] = 5'b00000; w[146][32] = 5'b10000; w[146][33] = 5'b00000; w[146][34] = 5'b01111; w[146][35] = 5'b01111; w[146][36] = 5'b01111; w[146][37] = 5'b10000; w[146][38] = 5'b00000; w[146][39] = 5'b01111; w[146][40] = 5'b00000; w[146][41] = 5'b00000; w[146][42] = 5'b00000; w[146][43] = 5'b00000; w[146][44] = 5'b01111; w[146][45] = 5'b10000; w[146][46] = 5'b10000; w[146][47] = 5'b00000; w[146][48] = 5'b01111; w[146][49] = 5'b01111; w[146][50] = 5'b01111; w[146][51] = 5'b10000; w[146][52] = 5'b10000; w[146][53] = 5'b01111; w[146][54] = 5'b00000; w[146][55] = 5'b00000; w[146][56] = 5'b00000; w[146][57] = 5'b00000; w[146][58] = 5'b10000; w[146][59] = 5'b10000; w[146][60] = 5'b10000; w[146][61] = 5'b10000; w[146][62] = 5'b01111; w[146][63] = 5'b01111; w[146][64] = 5'b00000; w[146][65] = 5'b10000; w[146][66] = 5'b10000; w[146][67] = 5'b10000; w[146][68] = 5'b00000; w[146][69] = 5'b00000; w[146][70] = 5'b00000; w[146][71] = 5'b00000; w[146][72] = 5'b10000; w[146][73] = 5'b10000; w[146][74] = 5'b10000; w[146][75] = 5'b10000; w[146][76] = 5'b01111; w[146][77] = 5'b01111; w[146][78] = 5'b00000; w[146][79] = 5'b10000; w[146][80] = 5'b10000; w[146][81] = 5'b10000; w[146][82] = 5'b00000; w[146][83] = 5'b00000; w[146][84] = 5'b00000; w[146][85] = 5'b00000; w[146][86] = 5'b10000; w[146][87] = 5'b10000; w[146][88] = 5'b10000; w[146][89] = 5'b10000; w[146][90] = 5'b01111; w[146][91] = 5'b01111; w[146][92] = 5'b00000; w[146][93] = 5'b10000; w[146][94] = 5'b10000; w[146][95] = 5'b00000; w[146][96] = 5'b00000; w[146][97] = 5'b00000; w[146][98] = 5'b00000; w[146][99] = 5'b00000; w[146][100] = 5'b10000; w[146][101] = 5'b10000; w[146][102] = 5'b10000; w[146][103] = 5'b00000; w[146][104] = 5'b01111; w[146][105] = 5'b01111; w[146][106] = 5'b10000; w[146][107] = 5'b10000; w[146][108] = 5'b10000; w[146][109] = 5'b10000; w[146][110] = 5'b00000; w[146][111] = 5'b00000; w[146][112] = 5'b00000; w[146][113] = 5'b00000; w[146][114] = 5'b10000; w[146][115] = 5'b10000; w[146][116] = 5'b10000; w[146][117] = 5'b00000; w[146][118] = 5'b01111; w[146][119] = 5'b01111; w[146][120] = 5'b10000; w[146][121] = 5'b10000; w[146][122] = 5'b10000; w[146][123] = 5'b10000; w[146][124] = 5'b00000; w[146][125] = 5'b00000; w[146][126] = 5'b00000; w[146][127] = 5'b00000; w[146][128] = 5'b10000; w[146][129] = 5'b10000; w[146][130] = 5'b10000; w[146][131] = 5'b00000; w[146][132] = 5'b01111; w[146][133] = 5'b01111; w[146][134] = 5'b10000; w[146][135] = 5'b10000; w[146][136] = 5'b10000; w[146][137] = 5'b10000; w[146][138] = 5'b00000; w[146][139] = 5'b00000; w[146][140] = 5'b00000; w[146][141] = 5'b00000; w[146][142] = 5'b10000; w[146][143] = 5'b10000; w[146][144] = 5'b10000; w[146][145] = 5'b00000; w[146][146] = 5'b00000; w[146][147] = 5'b01111; w[146][148] = 5'b10000; w[146][149] = 5'b10000; w[146][150] = 5'b10000; w[146][151] = 5'b10000; w[146][152] = 5'b00000; w[146][153] = 5'b00000; w[146][154] = 5'b00000; w[146][155] = 5'b00000; w[146][156] = 5'b00000; w[146][157] = 5'b10000; w[146][158] = 5'b10000; w[146][159] = 5'b00000; w[146][160] = 5'b01111; w[146][161] = 5'b01111; w[146][162] = 5'b10000; w[146][163] = 5'b10000; w[146][164] = 5'b10000; w[146][165] = 5'b00000; w[146][166] = 5'b00000; w[146][167] = 5'b00000; w[146][168] = 5'b00000; w[146][169] = 5'b00000; w[146][170] = 5'b00000; w[146][171] = 5'b10000; w[146][172] = 5'b10000; w[146][173] = 5'b00000; w[146][174] = 5'b01111; w[146][175] = 5'b01111; w[146][176] = 5'b10000; w[146][177] = 5'b10000; w[146][178] = 5'b10000; w[146][179] = 5'b00000; w[146][180] = 5'b00000; w[146][181] = 5'b00000; w[146][182] = 5'b00000; w[146][183] = 5'b00000; w[146][184] = 5'b00000; w[146][185] = 5'b00000; w[146][186] = 5'b00000; w[146][187] = 5'b00000; w[146][188] = 5'b00000; w[146][189] = 5'b00000; w[146][190] = 5'b00000; w[146][191] = 5'b00000; w[146][192] = 5'b00000; w[146][193] = 5'b00000; w[146][194] = 5'b00000; w[146][195] = 5'b00000; w[146][196] = 5'b00000; w[146][197] = 5'b00000; w[146][198] = 5'b00000; w[146][199] = 5'b00000; w[146][200] = 5'b00000; w[146][201] = 5'b00000; w[146][202] = 5'b00000; w[146][203] = 5'b00000; w[146][204] = 5'b00000; w[146][205] = 5'b00000; w[146][206] = 5'b00000; w[146][207] = 5'b00000; w[146][208] = 5'b00000; w[146][209] = 5'b00000; 
w[147][0] = 5'b10000; w[147][1] = 5'b10000; w[147][2] = 5'b10000; w[147][3] = 5'b10000; w[147][4] = 5'b10000; w[147][5] = 5'b10000; w[147][6] = 5'b10000; w[147][7] = 5'b10000; w[147][8] = 5'b10000; w[147][9] = 5'b10000; w[147][10] = 5'b10000; w[147][11] = 5'b10000; w[147][12] = 5'b10000; w[147][13] = 5'b10000; w[147][14] = 5'b10000; w[147][15] = 5'b10000; w[147][16] = 5'b10000; w[147][17] = 5'b10000; w[147][18] = 5'b10000; w[147][19] = 5'b10000; w[147][20] = 5'b10000; w[147][21] = 5'b10000; w[147][22] = 5'b10000; w[147][23] = 5'b10000; w[147][24] = 5'b10000; w[147][25] = 5'b10000; w[147][26] = 5'b10000; w[147][27] = 5'b10000; w[147][28] = 5'b10000; w[147][29] = 5'b10000; w[147][30] = 5'b00000; w[147][31] = 5'b01111; w[147][32] = 5'b00000; w[147][33] = 5'b01111; w[147][34] = 5'b00000; w[147][35] = 5'b00000; w[147][36] = 5'b00000; w[147][37] = 5'b00000; w[147][38] = 5'b01111; w[147][39] = 5'b00000; w[147][40] = 5'b10000; w[147][41] = 5'b10000; w[147][42] = 5'b10000; w[147][43] = 5'b10000; w[147][44] = 5'b00000; w[147][45] = 5'b00000; w[147][46] = 5'b00000; w[147][47] = 5'b01111; w[147][48] = 5'b00000; w[147][49] = 5'b00000; w[147][50] = 5'b00000; w[147][51] = 5'b00000; w[147][52] = 5'b00000; w[147][53] = 5'b00000; w[147][54] = 5'b10000; w[147][55] = 5'b10000; w[147][56] = 5'b10000; w[147][57] = 5'b10000; w[147][58] = 5'b10000; w[147][59] = 5'b10000; w[147][60] = 5'b10000; w[147][61] = 5'b00000; w[147][62] = 5'b01111; w[147][63] = 5'b01111; w[147][64] = 5'b10000; w[147][65] = 5'b10000; w[147][66] = 5'b10000; w[147][67] = 5'b10000; w[147][68] = 5'b10000; w[147][69] = 5'b10000; w[147][70] = 5'b10000; w[147][71] = 5'b10000; w[147][72] = 5'b10000; w[147][73] = 5'b10000; w[147][74] = 5'b00000; w[147][75] = 5'b00000; w[147][76] = 5'b01111; w[147][77] = 5'b01111; w[147][78] = 5'b10000; w[147][79] = 5'b00000; w[147][80] = 5'b10000; w[147][81] = 5'b10000; w[147][82] = 5'b10000; w[147][83] = 5'b10000; w[147][84] = 5'b10000; w[147][85] = 5'b10000; w[147][86] = 5'b10000; w[147][87] = 5'b10000; w[147][88] = 5'b00000; w[147][89] = 5'b00000; w[147][90] = 5'b01111; w[147][91] = 5'b01111; w[147][92] = 5'b10000; w[147][93] = 5'b00000; w[147][94] = 5'b00000; w[147][95] = 5'b10000; w[147][96] = 5'b10000; w[147][97] = 5'b10000; w[147][98] = 5'b10000; w[147][99] = 5'b10000; w[147][100] = 5'b10000; w[147][101] = 5'b10000; w[147][102] = 5'b00000; w[147][103] = 5'b10000; w[147][104] = 5'b01111; w[147][105] = 5'b01111; w[147][106] = 5'b10000; w[147][107] = 5'b10000; w[147][108] = 5'b10000; w[147][109] = 5'b10000; w[147][110] = 5'b10000; w[147][111] = 5'b10000; w[147][112] = 5'b10000; w[147][113] = 5'b10000; w[147][114] = 5'b10000; w[147][115] = 5'b10000; w[147][116] = 5'b00000; w[147][117] = 5'b10000; w[147][118] = 5'b01111; w[147][119] = 5'b01111; w[147][120] = 5'b10000; w[147][121] = 5'b10000; w[147][122] = 5'b10000; w[147][123] = 5'b10000; w[147][124] = 5'b10000; w[147][125] = 5'b10000; w[147][126] = 5'b10000; w[147][127] = 5'b10000; w[147][128] = 5'b10000; w[147][129] = 5'b10000; w[147][130] = 5'b00000; w[147][131] = 5'b10000; w[147][132] = 5'b01111; w[147][133] = 5'b01111; w[147][134] = 5'b00000; w[147][135] = 5'b00000; w[147][136] = 5'b10000; w[147][137] = 5'b10000; w[147][138] = 5'b10000; w[147][139] = 5'b10000; w[147][140] = 5'b10000; w[147][141] = 5'b10000; w[147][142] = 5'b10000; w[147][143] = 5'b10000; w[147][144] = 5'b10000; w[147][145] = 5'b10000; w[147][146] = 5'b01111; w[147][147] = 5'b00000; w[147][148] = 5'b00000; w[147][149] = 5'b10000; w[147][150] = 5'b10000; w[147][151] = 5'b10000; w[147][152] = 5'b10000; w[147][153] = 5'b10000; w[147][154] = 5'b10000; w[147][155] = 5'b10000; w[147][156] = 5'b10000; w[147][157] = 5'b10000; w[147][158] = 5'b10000; w[147][159] = 5'b10000; w[147][160] = 5'b00000; w[147][161] = 5'b00000; w[147][162] = 5'b00000; w[147][163] = 5'b10000; w[147][164] = 5'b10000; w[147][165] = 5'b10000; w[147][166] = 5'b10000; w[147][167] = 5'b10000; w[147][168] = 5'b10000; w[147][169] = 5'b10000; w[147][170] = 5'b10000; w[147][171] = 5'b00000; w[147][172] = 5'b10000; w[147][173] = 5'b10000; w[147][174] = 5'b00000; w[147][175] = 5'b00000; w[147][176] = 5'b00000; w[147][177] = 5'b10000; w[147][178] = 5'b00000; w[147][179] = 5'b10000; w[147][180] = 5'b10000; w[147][181] = 5'b10000; w[147][182] = 5'b10000; w[147][183] = 5'b10000; w[147][184] = 5'b10000; w[147][185] = 5'b10000; w[147][186] = 5'b10000; w[147][187] = 5'b10000; w[147][188] = 5'b10000; w[147][189] = 5'b10000; w[147][190] = 5'b10000; w[147][191] = 5'b10000; w[147][192] = 5'b10000; w[147][193] = 5'b10000; w[147][194] = 5'b10000; w[147][195] = 5'b10000; w[147][196] = 5'b10000; w[147][197] = 5'b10000; w[147][198] = 5'b10000; w[147][199] = 5'b10000; w[147][200] = 5'b10000; w[147][201] = 5'b10000; w[147][202] = 5'b10000; w[147][203] = 5'b10000; w[147][204] = 5'b10000; w[147][205] = 5'b10000; w[147][206] = 5'b10000; w[147][207] = 5'b10000; w[147][208] = 5'b10000; w[147][209] = 5'b10000; 
w[148][0] = 5'b01111; w[148][1] = 5'b01111; w[148][2] = 5'b01111; w[148][3] = 5'b01111; w[148][4] = 5'b01111; w[148][5] = 5'b01111; w[148][6] = 5'b01111; w[148][7] = 5'b01111; w[148][8] = 5'b01111; w[148][9] = 5'b01111; w[148][10] = 5'b01111; w[148][11] = 5'b01111; w[148][12] = 5'b01111; w[148][13] = 5'b01111; w[148][14] = 5'b01111; w[148][15] = 5'b01111; w[148][16] = 5'b01111; w[148][17] = 5'b01111; w[148][18] = 5'b01111; w[148][19] = 5'b01111; w[148][20] = 5'b01111; w[148][21] = 5'b01111; w[148][22] = 5'b01111; w[148][23] = 5'b01111; w[148][24] = 5'b01111; w[148][25] = 5'b01111; w[148][26] = 5'b01111; w[148][27] = 5'b01111; w[148][28] = 5'b01111; w[148][29] = 5'b01111; w[148][30] = 5'b00000; w[148][31] = 5'b01111; w[148][32] = 5'b00000; w[148][33] = 5'b10000; w[148][34] = 5'b10000; w[148][35] = 5'b10000; w[148][36] = 5'b10000; w[148][37] = 5'b00000; w[148][38] = 5'b01111; w[148][39] = 5'b00000; w[148][40] = 5'b01111; w[148][41] = 5'b01111; w[148][42] = 5'b01111; w[148][43] = 5'b01111; w[148][44] = 5'b00000; w[148][45] = 5'b00000; w[148][46] = 5'b00000; w[148][47] = 5'b10000; w[148][48] = 5'b10000; w[148][49] = 5'b10000; w[148][50] = 5'b10000; w[148][51] = 5'b00000; w[148][52] = 5'b00000; w[148][53] = 5'b00000; w[148][54] = 5'b01111; w[148][55] = 5'b01111; w[148][56] = 5'b01111; w[148][57] = 5'b01111; w[148][58] = 5'b00000; w[148][59] = 5'b01111; w[148][60] = 5'b01111; w[148][61] = 5'b01111; w[148][62] = 5'b00000; w[148][63] = 5'b10000; w[148][64] = 5'b01111; w[148][65] = 5'b01111; w[148][66] = 5'b01111; w[148][67] = 5'b00000; w[148][68] = 5'b01111; w[148][69] = 5'b01111; w[148][70] = 5'b01111; w[148][71] = 5'b01111; w[148][72] = 5'b00000; w[148][73] = 5'b01111; w[148][74] = 5'b01111; w[148][75] = 5'b01111; w[148][76] = 5'b00000; w[148][77] = 5'b10000; w[148][78] = 5'b01111; w[148][79] = 5'b01111; w[148][80] = 5'b01111; w[148][81] = 5'b00000; w[148][82] = 5'b01111; w[148][83] = 5'b01111; w[148][84] = 5'b01111; w[148][85] = 5'b01111; w[148][86] = 5'b00000; w[148][87] = 5'b01111; w[148][88] = 5'b01111; w[148][89] = 5'b01111; w[148][90] = 5'b00000; w[148][91] = 5'b00000; w[148][92] = 5'b01111; w[148][93] = 5'b01111; w[148][94] = 5'b01111; w[148][95] = 5'b01111; w[148][96] = 5'b01111; w[148][97] = 5'b01111; w[148][98] = 5'b01111; w[148][99] = 5'b01111; w[148][100] = 5'b00000; w[148][101] = 5'b01111; w[148][102] = 5'b01111; w[148][103] = 5'b01111; w[148][104] = 5'b00000; w[148][105] = 5'b00000; w[148][106] = 5'b00000; w[148][107] = 5'b01111; w[148][108] = 5'b01111; w[148][109] = 5'b00000; w[148][110] = 5'b01111; w[148][111] = 5'b01111; w[148][112] = 5'b01111; w[148][113] = 5'b01111; w[148][114] = 5'b00000; w[148][115] = 5'b01111; w[148][116] = 5'b01111; w[148][117] = 5'b01111; w[148][118] = 5'b00000; w[148][119] = 5'b00000; w[148][120] = 5'b01111; w[148][121] = 5'b01111; w[148][122] = 5'b01111; w[148][123] = 5'b00000; w[148][124] = 5'b01111; w[148][125] = 5'b01111; w[148][126] = 5'b01111; w[148][127] = 5'b01111; w[148][128] = 5'b00000; w[148][129] = 5'b01111; w[148][130] = 5'b01111; w[148][131] = 5'b01111; w[148][132] = 5'b10000; w[148][133] = 5'b00000; w[148][134] = 5'b01111; w[148][135] = 5'b01111; w[148][136] = 5'b01111; w[148][137] = 5'b00000; w[148][138] = 5'b01111; w[148][139] = 5'b01111; w[148][140] = 5'b01111; w[148][141] = 5'b01111; w[148][142] = 5'b00000; w[148][143] = 5'b01111; w[148][144] = 5'b01111; w[148][145] = 5'b01111; w[148][146] = 5'b10000; w[148][147] = 5'b00000; w[148][148] = 5'b00000; w[148][149] = 5'b01111; w[148][150] = 5'b01111; w[148][151] = 5'b00000; w[148][152] = 5'b01111; w[148][153] = 5'b01111; w[148][154] = 5'b01111; w[148][155] = 5'b01111; w[148][156] = 5'b01111; w[148][157] = 5'b01111; w[148][158] = 5'b01111; w[148][159] = 5'b10000; w[148][160] = 5'b10000; w[148][161] = 5'b10000; w[148][162] = 5'b00000; w[148][163] = 5'b01111; w[148][164] = 5'b01111; w[148][165] = 5'b01111; w[148][166] = 5'b01111; w[148][167] = 5'b01111; w[148][168] = 5'b01111; w[148][169] = 5'b01111; w[148][170] = 5'b01111; w[148][171] = 5'b01111; w[148][172] = 5'b01111; w[148][173] = 5'b10000; w[148][174] = 5'b10000; w[148][175] = 5'b10000; w[148][176] = 5'b00000; w[148][177] = 5'b01111; w[148][178] = 5'b01111; w[148][179] = 5'b01111; w[148][180] = 5'b01111; w[148][181] = 5'b01111; w[148][182] = 5'b01111; w[148][183] = 5'b01111; w[148][184] = 5'b01111; w[148][185] = 5'b01111; w[148][186] = 5'b01111; w[148][187] = 5'b01111; w[148][188] = 5'b01111; w[148][189] = 5'b01111; w[148][190] = 5'b01111; w[148][191] = 5'b01111; w[148][192] = 5'b01111; w[148][193] = 5'b01111; w[148][194] = 5'b01111; w[148][195] = 5'b01111; w[148][196] = 5'b01111; w[148][197] = 5'b01111; w[148][198] = 5'b01111; w[148][199] = 5'b01111; w[148][200] = 5'b01111; w[148][201] = 5'b01111; w[148][202] = 5'b01111; w[148][203] = 5'b01111; w[148][204] = 5'b01111; w[148][205] = 5'b01111; w[148][206] = 5'b01111; w[148][207] = 5'b01111; w[148][208] = 5'b01111; w[148][209] = 5'b01111; 
w[149][0] = 5'b00000; w[149][1] = 5'b00000; w[149][2] = 5'b00000; w[149][3] = 5'b00000; w[149][4] = 5'b00000; w[149][5] = 5'b00000; w[149][6] = 5'b00000; w[149][7] = 5'b00000; w[149][8] = 5'b00000; w[149][9] = 5'b00000; w[149][10] = 5'b00000; w[149][11] = 5'b00000; w[149][12] = 5'b00000; w[149][13] = 5'b00000; w[149][14] = 5'b00000; w[149][15] = 5'b00000; w[149][16] = 5'b00000; w[149][17] = 5'b00000; w[149][18] = 5'b00000; w[149][19] = 5'b00000; w[149][20] = 5'b00000; w[149][21] = 5'b00000; w[149][22] = 5'b00000; w[149][23] = 5'b00000; w[149][24] = 5'b00000; w[149][25] = 5'b00000; w[149][26] = 5'b00000; w[149][27] = 5'b00000; w[149][28] = 5'b00000; w[149][29] = 5'b00000; w[149][30] = 5'b10000; w[149][31] = 5'b00000; w[149][32] = 5'b01111; w[149][33] = 5'b00000; w[149][34] = 5'b10000; w[149][35] = 5'b10000; w[149][36] = 5'b10000; w[149][37] = 5'b01111; w[149][38] = 5'b00000; w[149][39] = 5'b10000; w[149][40] = 5'b00000; w[149][41] = 5'b00000; w[149][42] = 5'b00000; w[149][43] = 5'b00000; w[149][44] = 5'b10000; w[149][45] = 5'b01111; w[149][46] = 5'b01111; w[149][47] = 5'b00000; w[149][48] = 5'b10000; w[149][49] = 5'b10000; w[149][50] = 5'b10000; w[149][51] = 5'b01111; w[149][52] = 5'b01111; w[149][53] = 5'b10000; w[149][54] = 5'b00000; w[149][55] = 5'b00000; w[149][56] = 5'b00000; w[149][57] = 5'b00000; w[149][58] = 5'b01111; w[149][59] = 5'b01111; w[149][60] = 5'b01111; w[149][61] = 5'b01111; w[149][62] = 5'b10000; w[149][63] = 5'b10000; w[149][64] = 5'b00000; w[149][65] = 5'b01111; w[149][66] = 5'b01111; w[149][67] = 5'b01111; w[149][68] = 5'b00000; w[149][69] = 5'b00000; w[149][70] = 5'b00000; w[149][71] = 5'b00000; w[149][72] = 5'b01111; w[149][73] = 5'b01111; w[149][74] = 5'b01111; w[149][75] = 5'b01111; w[149][76] = 5'b10000; w[149][77] = 5'b10000; w[149][78] = 5'b00000; w[149][79] = 5'b01111; w[149][80] = 5'b01111; w[149][81] = 5'b01111; w[149][82] = 5'b00000; w[149][83] = 5'b00000; w[149][84] = 5'b00000; w[149][85] = 5'b00000; w[149][86] = 5'b01111; w[149][87] = 5'b01111; w[149][88] = 5'b01111; w[149][89] = 5'b01111; w[149][90] = 5'b10000; w[149][91] = 5'b10000; w[149][92] = 5'b00000; w[149][93] = 5'b01111; w[149][94] = 5'b01111; w[149][95] = 5'b00000; w[149][96] = 5'b00000; w[149][97] = 5'b00000; w[149][98] = 5'b00000; w[149][99] = 5'b00000; w[149][100] = 5'b01111; w[149][101] = 5'b01111; w[149][102] = 5'b01111; w[149][103] = 5'b00000; w[149][104] = 5'b10000; w[149][105] = 5'b10000; w[149][106] = 5'b01111; w[149][107] = 5'b01111; w[149][108] = 5'b01111; w[149][109] = 5'b01111; w[149][110] = 5'b00000; w[149][111] = 5'b00000; w[149][112] = 5'b00000; w[149][113] = 5'b00000; w[149][114] = 5'b01111; w[149][115] = 5'b01111; w[149][116] = 5'b01111; w[149][117] = 5'b00000; w[149][118] = 5'b10000; w[149][119] = 5'b10000; w[149][120] = 5'b01111; w[149][121] = 5'b01111; w[149][122] = 5'b01111; w[149][123] = 5'b01111; w[149][124] = 5'b00000; w[149][125] = 5'b00000; w[149][126] = 5'b00000; w[149][127] = 5'b00000; w[149][128] = 5'b01111; w[149][129] = 5'b01111; w[149][130] = 5'b01111; w[149][131] = 5'b00000; w[149][132] = 5'b10000; w[149][133] = 5'b10000; w[149][134] = 5'b01111; w[149][135] = 5'b01111; w[149][136] = 5'b01111; w[149][137] = 5'b01111; w[149][138] = 5'b00000; w[149][139] = 5'b00000; w[149][140] = 5'b00000; w[149][141] = 5'b00000; w[149][142] = 5'b01111; w[149][143] = 5'b01111; w[149][144] = 5'b01111; w[149][145] = 5'b00000; w[149][146] = 5'b10000; w[149][147] = 5'b10000; w[149][148] = 5'b01111; w[149][149] = 5'b00000; w[149][150] = 5'b01111; w[149][151] = 5'b01111; w[149][152] = 5'b00000; w[149][153] = 5'b00000; w[149][154] = 5'b00000; w[149][155] = 5'b00000; w[149][156] = 5'b00000; w[149][157] = 5'b01111; w[149][158] = 5'b01111; w[149][159] = 5'b00000; w[149][160] = 5'b10000; w[149][161] = 5'b10000; w[149][162] = 5'b01111; w[149][163] = 5'b01111; w[149][164] = 5'b01111; w[149][165] = 5'b00000; w[149][166] = 5'b00000; w[149][167] = 5'b00000; w[149][168] = 5'b00000; w[149][169] = 5'b00000; w[149][170] = 5'b00000; w[149][171] = 5'b01111; w[149][172] = 5'b01111; w[149][173] = 5'b00000; w[149][174] = 5'b10000; w[149][175] = 5'b10000; w[149][176] = 5'b01111; w[149][177] = 5'b01111; w[149][178] = 5'b01111; w[149][179] = 5'b00000; w[149][180] = 5'b00000; w[149][181] = 5'b00000; w[149][182] = 5'b00000; w[149][183] = 5'b00000; w[149][184] = 5'b00000; w[149][185] = 5'b00000; w[149][186] = 5'b00000; w[149][187] = 5'b00000; w[149][188] = 5'b00000; w[149][189] = 5'b00000; w[149][190] = 5'b00000; w[149][191] = 5'b00000; w[149][192] = 5'b00000; w[149][193] = 5'b00000; w[149][194] = 5'b00000; w[149][195] = 5'b00000; w[149][196] = 5'b00000; w[149][197] = 5'b00000; w[149][198] = 5'b00000; w[149][199] = 5'b00000; w[149][200] = 5'b00000; w[149][201] = 5'b00000; w[149][202] = 5'b00000; w[149][203] = 5'b00000; w[149][204] = 5'b00000; w[149][205] = 5'b00000; w[149][206] = 5'b00000; w[149][207] = 5'b00000; w[149][208] = 5'b00000; w[149][209] = 5'b00000; 
w[150][0] = 5'b00000; w[150][1] = 5'b00000; w[150][2] = 5'b00000; w[150][3] = 5'b00000; w[150][4] = 5'b00000; w[150][5] = 5'b00000; w[150][6] = 5'b00000; w[150][7] = 5'b00000; w[150][8] = 5'b00000; w[150][9] = 5'b00000; w[150][10] = 5'b00000; w[150][11] = 5'b00000; w[150][12] = 5'b00000; w[150][13] = 5'b00000; w[150][14] = 5'b00000; w[150][15] = 5'b00000; w[150][16] = 5'b00000; w[150][17] = 5'b00000; w[150][18] = 5'b00000; w[150][19] = 5'b00000; w[150][20] = 5'b00000; w[150][21] = 5'b00000; w[150][22] = 5'b00000; w[150][23] = 5'b00000; w[150][24] = 5'b00000; w[150][25] = 5'b00000; w[150][26] = 5'b00000; w[150][27] = 5'b00000; w[150][28] = 5'b00000; w[150][29] = 5'b00000; w[150][30] = 5'b10000; w[150][31] = 5'b00000; w[150][32] = 5'b01111; w[150][33] = 5'b00000; w[150][34] = 5'b10000; w[150][35] = 5'b10000; w[150][36] = 5'b10000; w[150][37] = 5'b01111; w[150][38] = 5'b00000; w[150][39] = 5'b10000; w[150][40] = 5'b00000; w[150][41] = 5'b00000; w[150][42] = 5'b00000; w[150][43] = 5'b00000; w[150][44] = 5'b10000; w[150][45] = 5'b01111; w[150][46] = 5'b01111; w[150][47] = 5'b00000; w[150][48] = 5'b10000; w[150][49] = 5'b10000; w[150][50] = 5'b10000; w[150][51] = 5'b01111; w[150][52] = 5'b01111; w[150][53] = 5'b10000; w[150][54] = 5'b00000; w[150][55] = 5'b00000; w[150][56] = 5'b00000; w[150][57] = 5'b00000; w[150][58] = 5'b01111; w[150][59] = 5'b01111; w[150][60] = 5'b01111; w[150][61] = 5'b01111; w[150][62] = 5'b10000; w[150][63] = 5'b10000; w[150][64] = 5'b00000; w[150][65] = 5'b01111; w[150][66] = 5'b01111; w[150][67] = 5'b01111; w[150][68] = 5'b00000; w[150][69] = 5'b00000; w[150][70] = 5'b00000; w[150][71] = 5'b00000; w[150][72] = 5'b01111; w[150][73] = 5'b01111; w[150][74] = 5'b01111; w[150][75] = 5'b01111; w[150][76] = 5'b10000; w[150][77] = 5'b10000; w[150][78] = 5'b00000; w[150][79] = 5'b01111; w[150][80] = 5'b01111; w[150][81] = 5'b01111; w[150][82] = 5'b00000; w[150][83] = 5'b00000; w[150][84] = 5'b00000; w[150][85] = 5'b00000; w[150][86] = 5'b01111; w[150][87] = 5'b01111; w[150][88] = 5'b01111; w[150][89] = 5'b01111; w[150][90] = 5'b10000; w[150][91] = 5'b10000; w[150][92] = 5'b00000; w[150][93] = 5'b01111; w[150][94] = 5'b01111; w[150][95] = 5'b00000; w[150][96] = 5'b00000; w[150][97] = 5'b00000; w[150][98] = 5'b00000; w[150][99] = 5'b00000; w[150][100] = 5'b01111; w[150][101] = 5'b01111; w[150][102] = 5'b01111; w[150][103] = 5'b00000; w[150][104] = 5'b10000; w[150][105] = 5'b10000; w[150][106] = 5'b01111; w[150][107] = 5'b01111; w[150][108] = 5'b01111; w[150][109] = 5'b01111; w[150][110] = 5'b00000; w[150][111] = 5'b00000; w[150][112] = 5'b00000; w[150][113] = 5'b00000; w[150][114] = 5'b01111; w[150][115] = 5'b01111; w[150][116] = 5'b01111; w[150][117] = 5'b00000; w[150][118] = 5'b10000; w[150][119] = 5'b10000; w[150][120] = 5'b01111; w[150][121] = 5'b01111; w[150][122] = 5'b01111; w[150][123] = 5'b01111; w[150][124] = 5'b00000; w[150][125] = 5'b00000; w[150][126] = 5'b00000; w[150][127] = 5'b00000; w[150][128] = 5'b01111; w[150][129] = 5'b01111; w[150][130] = 5'b01111; w[150][131] = 5'b00000; w[150][132] = 5'b10000; w[150][133] = 5'b10000; w[150][134] = 5'b01111; w[150][135] = 5'b01111; w[150][136] = 5'b01111; w[150][137] = 5'b01111; w[150][138] = 5'b00000; w[150][139] = 5'b00000; w[150][140] = 5'b00000; w[150][141] = 5'b00000; w[150][142] = 5'b01111; w[150][143] = 5'b01111; w[150][144] = 5'b01111; w[150][145] = 5'b00000; w[150][146] = 5'b10000; w[150][147] = 5'b10000; w[150][148] = 5'b01111; w[150][149] = 5'b01111; w[150][150] = 5'b00000; w[150][151] = 5'b01111; w[150][152] = 5'b00000; w[150][153] = 5'b00000; w[150][154] = 5'b00000; w[150][155] = 5'b00000; w[150][156] = 5'b00000; w[150][157] = 5'b01111; w[150][158] = 5'b01111; w[150][159] = 5'b00000; w[150][160] = 5'b10000; w[150][161] = 5'b10000; w[150][162] = 5'b01111; w[150][163] = 5'b01111; w[150][164] = 5'b01111; w[150][165] = 5'b00000; w[150][166] = 5'b00000; w[150][167] = 5'b00000; w[150][168] = 5'b00000; w[150][169] = 5'b00000; w[150][170] = 5'b00000; w[150][171] = 5'b01111; w[150][172] = 5'b01111; w[150][173] = 5'b00000; w[150][174] = 5'b10000; w[150][175] = 5'b10000; w[150][176] = 5'b01111; w[150][177] = 5'b01111; w[150][178] = 5'b01111; w[150][179] = 5'b00000; w[150][180] = 5'b00000; w[150][181] = 5'b00000; w[150][182] = 5'b00000; w[150][183] = 5'b00000; w[150][184] = 5'b00000; w[150][185] = 5'b00000; w[150][186] = 5'b00000; w[150][187] = 5'b00000; w[150][188] = 5'b00000; w[150][189] = 5'b00000; w[150][190] = 5'b00000; w[150][191] = 5'b00000; w[150][192] = 5'b00000; w[150][193] = 5'b00000; w[150][194] = 5'b00000; w[150][195] = 5'b00000; w[150][196] = 5'b00000; w[150][197] = 5'b00000; w[150][198] = 5'b00000; w[150][199] = 5'b00000; w[150][200] = 5'b00000; w[150][201] = 5'b00000; w[150][202] = 5'b00000; w[150][203] = 5'b00000; w[150][204] = 5'b00000; w[150][205] = 5'b00000; w[150][206] = 5'b00000; w[150][207] = 5'b00000; w[150][208] = 5'b00000; w[150][209] = 5'b00000; 
w[151][0] = 5'b01111; w[151][1] = 5'b01111; w[151][2] = 5'b01111; w[151][3] = 5'b01111; w[151][4] = 5'b01111; w[151][5] = 5'b01111; w[151][6] = 5'b01111; w[151][7] = 5'b01111; w[151][8] = 5'b01111; w[151][9] = 5'b01111; w[151][10] = 5'b01111; w[151][11] = 5'b01111; w[151][12] = 5'b01111; w[151][13] = 5'b01111; w[151][14] = 5'b01111; w[151][15] = 5'b01111; w[151][16] = 5'b01111; w[151][17] = 5'b01111; w[151][18] = 5'b01111; w[151][19] = 5'b01111; w[151][20] = 5'b01111; w[151][21] = 5'b01111; w[151][22] = 5'b01111; w[151][23] = 5'b01111; w[151][24] = 5'b01111; w[151][25] = 5'b01111; w[151][26] = 5'b01111; w[151][27] = 5'b01111; w[151][28] = 5'b01111; w[151][29] = 5'b01111; w[151][30] = 5'b00000; w[151][31] = 5'b10000; w[151][32] = 5'b00000; w[151][33] = 5'b10000; w[151][34] = 5'b00000; w[151][35] = 5'b00000; w[151][36] = 5'b00000; w[151][37] = 5'b00000; w[151][38] = 5'b10000; w[151][39] = 5'b00000; w[151][40] = 5'b01111; w[151][41] = 5'b01111; w[151][42] = 5'b01111; w[151][43] = 5'b01111; w[151][44] = 5'b00000; w[151][45] = 5'b00000; w[151][46] = 5'b00000; w[151][47] = 5'b10000; w[151][48] = 5'b00000; w[151][49] = 5'b00000; w[151][50] = 5'b00000; w[151][51] = 5'b00000; w[151][52] = 5'b00000; w[151][53] = 5'b00000; w[151][54] = 5'b01111; w[151][55] = 5'b01111; w[151][56] = 5'b01111; w[151][57] = 5'b01111; w[151][58] = 5'b01111; w[151][59] = 5'b01111; w[151][60] = 5'b01111; w[151][61] = 5'b00000; w[151][62] = 5'b10000; w[151][63] = 5'b10000; w[151][64] = 5'b01111; w[151][65] = 5'b01111; w[151][66] = 5'b01111; w[151][67] = 5'b01111; w[151][68] = 5'b01111; w[151][69] = 5'b01111; w[151][70] = 5'b01111; w[151][71] = 5'b01111; w[151][72] = 5'b01111; w[151][73] = 5'b01111; w[151][74] = 5'b00000; w[151][75] = 5'b00000; w[151][76] = 5'b10000; w[151][77] = 5'b10000; w[151][78] = 5'b01111; w[151][79] = 5'b00000; w[151][80] = 5'b01111; w[151][81] = 5'b01111; w[151][82] = 5'b01111; w[151][83] = 5'b01111; w[151][84] = 5'b01111; w[151][85] = 5'b01111; w[151][86] = 5'b01111; w[151][87] = 5'b01111; w[151][88] = 5'b00000; w[151][89] = 5'b00000; w[151][90] = 5'b10000; w[151][91] = 5'b10000; w[151][92] = 5'b01111; w[151][93] = 5'b00000; w[151][94] = 5'b00000; w[151][95] = 5'b01111; w[151][96] = 5'b01111; w[151][97] = 5'b01111; w[151][98] = 5'b01111; w[151][99] = 5'b01111; w[151][100] = 5'b01111; w[151][101] = 5'b01111; w[151][102] = 5'b00000; w[151][103] = 5'b01111; w[151][104] = 5'b10000; w[151][105] = 5'b10000; w[151][106] = 5'b01111; w[151][107] = 5'b01111; w[151][108] = 5'b01111; w[151][109] = 5'b01111; w[151][110] = 5'b01111; w[151][111] = 5'b01111; w[151][112] = 5'b01111; w[151][113] = 5'b01111; w[151][114] = 5'b01111; w[151][115] = 5'b01111; w[151][116] = 5'b00000; w[151][117] = 5'b01111; w[151][118] = 5'b10000; w[151][119] = 5'b10000; w[151][120] = 5'b01111; w[151][121] = 5'b01111; w[151][122] = 5'b01111; w[151][123] = 5'b01111; w[151][124] = 5'b01111; w[151][125] = 5'b01111; w[151][126] = 5'b01111; w[151][127] = 5'b01111; w[151][128] = 5'b01111; w[151][129] = 5'b01111; w[151][130] = 5'b00000; w[151][131] = 5'b01111; w[151][132] = 5'b10000; w[151][133] = 5'b10000; w[151][134] = 5'b00000; w[151][135] = 5'b00000; w[151][136] = 5'b01111; w[151][137] = 5'b01111; w[151][138] = 5'b01111; w[151][139] = 5'b01111; w[151][140] = 5'b01111; w[151][141] = 5'b01111; w[151][142] = 5'b01111; w[151][143] = 5'b01111; w[151][144] = 5'b01111; w[151][145] = 5'b01111; w[151][146] = 5'b10000; w[151][147] = 5'b10000; w[151][148] = 5'b00000; w[151][149] = 5'b01111; w[151][150] = 5'b01111; w[151][151] = 5'b00000; w[151][152] = 5'b01111; w[151][153] = 5'b01111; w[151][154] = 5'b01111; w[151][155] = 5'b01111; w[151][156] = 5'b01111; w[151][157] = 5'b01111; w[151][158] = 5'b01111; w[151][159] = 5'b01111; w[151][160] = 5'b00000; w[151][161] = 5'b00000; w[151][162] = 5'b00000; w[151][163] = 5'b01111; w[151][164] = 5'b01111; w[151][165] = 5'b01111; w[151][166] = 5'b01111; w[151][167] = 5'b01111; w[151][168] = 5'b01111; w[151][169] = 5'b01111; w[151][170] = 5'b01111; w[151][171] = 5'b00000; w[151][172] = 5'b01111; w[151][173] = 5'b01111; w[151][174] = 5'b00000; w[151][175] = 5'b00000; w[151][176] = 5'b00000; w[151][177] = 5'b01111; w[151][178] = 5'b00000; w[151][179] = 5'b01111; w[151][180] = 5'b01111; w[151][181] = 5'b01111; w[151][182] = 5'b01111; w[151][183] = 5'b01111; w[151][184] = 5'b01111; w[151][185] = 5'b01111; w[151][186] = 5'b01111; w[151][187] = 5'b01111; w[151][188] = 5'b01111; w[151][189] = 5'b01111; w[151][190] = 5'b01111; w[151][191] = 5'b01111; w[151][192] = 5'b01111; w[151][193] = 5'b01111; w[151][194] = 5'b01111; w[151][195] = 5'b01111; w[151][196] = 5'b01111; w[151][197] = 5'b01111; w[151][198] = 5'b01111; w[151][199] = 5'b01111; w[151][200] = 5'b01111; w[151][201] = 5'b01111; w[151][202] = 5'b01111; w[151][203] = 5'b01111; w[151][204] = 5'b01111; w[151][205] = 5'b01111; w[151][206] = 5'b01111; w[151][207] = 5'b01111; w[151][208] = 5'b01111; w[151][209] = 5'b01111; 
w[152][0] = 5'b01111; w[152][1] = 5'b01111; w[152][2] = 5'b01111; w[152][3] = 5'b01111; w[152][4] = 5'b01111; w[152][5] = 5'b01111; w[152][6] = 5'b01111; w[152][7] = 5'b01111; w[152][8] = 5'b01111; w[152][9] = 5'b01111; w[152][10] = 5'b01111; w[152][11] = 5'b01111; w[152][12] = 5'b01111; w[152][13] = 5'b01111; w[152][14] = 5'b01111; w[152][15] = 5'b01111; w[152][16] = 5'b01111; w[152][17] = 5'b01111; w[152][18] = 5'b01111; w[152][19] = 5'b01111; w[152][20] = 5'b01111; w[152][21] = 5'b01111; w[152][22] = 5'b01111; w[152][23] = 5'b01111; w[152][24] = 5'b01111; w[152][25] = 5'b01111; w[152][26] = 5'b01111; w[152][27] = 5'b01111; w[152][28] = 5'b01111; w[152][29] = 5'b01111; w[152][30] = 5'b01111; w[152][31] = 5'b00000; w[152][32] = 5'b10000; w[152][33] = 5'b10000; w[152][34] = 5'b10000; w[152][35] = 5'b10000; w[152][36] = 5'b10000; w[152][37] = 5'b10000; w[152][38] = 5'b00000; w[152][39] = 5'b01111; w[152][40] = 5'b01111; w[152][41] = 5'b01111; w[152][42] = 5'b01111; w[152][43] = 5'b01111; w[152][44] = 5'b01111; w[152][45] = 5'b10000; w[152][46] = 5'b10000; w[152][47] = 5'b10000; w[152][48] = 5'b10000; w[152][49] = 5'b10000; w[152][50] = 5'b10000; w[152][51] = 5'b10000; w[152][52] = 5'b10000; w[152][53] = 5'b01111; w[152][54] = 5'b01111; w[152][55] = 5'b01111; w[152][56] = 5'b01111; w[152][57] = 5'b01111; w[152][58] = 5'b01111; w[152][59] = 5'b00000; w[152][60] = 5'b00000; w[152][61] = 5'b01111; w[152][62] = 5'b10000; w[152][63] = 5'b00000; w[152][64] = 5'b01111; w[152][65] = 5'b00000; w[152][66] = 5'b00000; w[152][67] = 5'b01111; w[152][68] = 5'b01111; w[152][69] = 5'b01111; w[152][70] = 5'b01111; w[152][71] = 5'b01111; w[152][72] = 5'b01111; w[152][73] = 5'b00000; w[152][74] = 5'b01111; w[152][75] = 5'b01111; w[152][76] = 5'b10000; w[152][77] = 5'b00000; w[152][78] = 5'b01111; w[152][79] = 5'b01111; w[152][80] = 5'b00000; w[152][81] = 5'b01111; w[152][82] = 5'b01111; w[152][83] = 5'b01111; w[152][84] = 5'b01111; w[152][85] = 5'b01111; w[152][86] = 5'b01111; w[152][87] = 5'b00000; w[152][88] = 5'b01111; w[152][89] = 5'b01111; w[152][90] = 5'b10000; w[152][91] = 5'b10000; w[152][92] = 5'b01111; w[152][93] = 5'b01111; w[152][94] = 5'b01111; w[152][95] = 5'b01111; w[152][96] = 5'b01111; w[152][97] = 5'b01111; w[152][98] = 5'b01111; w[152][99] = 5'b01111; w[152][100] = 5'b01111; w[152][101] = 5'b00000; w[152][102] = 5'b01111; w[152][103] = 5'b01111; w[152][104] = 5'b10000; w[152][105] = 5'b10000; w[152][106] = 5'b01111; w[152][107] = 5'b00000; w[152][108] = 5'b00000; w[152][109] = 5'b01111; w[152][110] = 5'b01111; w[152][111] = 5'b01111; w[152][112] = 5'b01111; w[152][113] = 5'b01111; w[152][114] = 5'b01111; w[152][115] = 5'b00000; w[152][116] = 5'b01111; w[152][117] = 5'b01111; w[152][118] = 5'b10000; w[152][119] = 5'b10000; w[152][120] = 5'b00000; w[152][121] = 5'b00000; w[152][122] = 5'b00000; w[152][123] = 5'b01111; w[152][124] = 5'b01111; w[152][125] = 5'b01111; w[152][126] = 5'b01111; w[152][127] = 5'b01111; w[152][128] = 5'b01111; w[152][129] = 5'b00000; w[152][130] = 5'b01111; w[152][131] = 5'b01111; w[152][132] = 5'b00000; w[152][133] = 5'b10000; w[152][134] = 5'b01111; w[152][135] = 5'b01111; w[152][136] = 5'b00000; w[152][137] = 5'b01111; w[152][138] = 5'b01111; w[152][139] = 5'b01111; w[152][140] = 5'b01111; w[152][141] = 5'b01111; w[152][142] = 5'b01111; w[152][143] = 5'b00000; w[152][144] = 5'b00000; w[152][145] = 5'b01111; w[152][146] = 5'b00000; w[152][147] = 5'b10000; w[152][148] = 5'b01111; w[152][149] = 5'b00000; w[152][150] = 5'b00000; w[152][151] = 5'b01111; w[152][152] = 5'b00000; w[152][153] = 5'b01111; w[152][154] = 5'b01111; w[152][155] = 5'b01111; w[152][156] = 5'b01111; w[152][157] = 5'b00000; w[152][158] = 5'b00000; w[152][159] = 5'b00000; w[152][160] = 5'b10000; w[152][161] = 5'b10000; w[152][162] = 5'b10000; w[152][163] = 5'b00000; w[152][164] = 5'b00000; w[152][165] = 5'b01111; w[152][166] = 5'b01111; w[152][167] = 5'b01111; w[152][168] = 5'b01111; w[152][169] = 5'b01111; w[152][170] = 5'b01111; w[152][171] = 5'b01111; w[152][172] = 5'b00000; w[152][173] = 5'b00000; w[152][174] = 5'b10000; w[152][175] = 5'b10000; w[152][176] = 5'b10000; w[152][177] = 5'b00000; w[152][178] = 5'b01111; w[152][179] = 5'b01111; w[152][180] = 5'b01111; w[152][181] = 5'b01111; w[152][182] = 5'b01111; w[152][183] = 5'b01111; w[152][184] = 5'b01111; w[152][185] = 5'b01111; w[152][186] = 5'b01111; w[152][187] = 5'b01111; w[152][188] = 5'b01111; w[152][189] = 5'b01111; w[152][190] = 5'b01111; w[152][191] = 5'b01111; w[152][192] = 5'b01111; w[152][193] = 5'b01111; w[152][194] = 5'b01111; w[152][195] = 5'b01111; w[152][196] = 5'b01111; w[152][197] = 5'b01111; w[152][198] = 5'b01111; w[152][199] = 5'b01111; w[152][200] = 5'b01111; w[152][201] = 5'b01111; w[152][202] = 5'b01111; w[152][203] = 5'b01111; w[152][204] = 5'b01111; w[152][205] = 5'b01111; w[152][206] = 5'b01111; w[152][207] = 5'b01111; w[152][208] = 5'b01111; w[152][209] = 5'b01111; 
w[153][0] = 5'b01111; w[153][1] = 5'b01111; w[153][2] = 5'b01111; w[153][3] = 5'b01111; w[153][4] = 5'b01111; w[153][5] = 5'b01111; w[153][6] = 5'b01111; w[153][7] = 5'b01111; w[153][8] = 5'b01111; w[153][9] = 5'b01111; w[153][10] = 5'b01111; w[153][11] = 5'b01111; w[153][12] = 5'b01111; w[153][13] = 5'b01111; w[153][14] = 5'b01111; w[153][15] = 5'b01111; w[153][16] = 5'b01111; w[153][17] = 5'b01111; w[153][18] = 5'b01111; w[153][19] = 5'b01111; w[153][20] = 5'b01111; w[153][21] = 5'b01111; w[153][22] = 5'b01111; w[153][23] = 5'b01111; w[153][24] = 5'b01111; w[153][25] = 5'b01111; w[153][26] = 5'b01111; w[153][27] = 5'b01111; w[153][28] = 5'b01111; w[153][29] = 5'b01111; w[153][30] = 5'b01111; w[153][31] = 5'b00000; w[153][32] = 5'b10000; w[153][33] = 5'b10000; w[153][34] = 5'b10000; w[153][35] = 5'b10000; w[153][36] = 5'b10000; w[153][37] = 5'b10000; w[153][38] = 5'b00000; w[153][39] = 5'b01111; w[153][40] = 5'b01111; w[153][41] = 5'b01111; w[153][42] = 5'b01111; w[153][43] = 5'b01111; w[153][44] = 5'b01111; w[153][45] = 5'b10000; w[153][46] = 5'b10000; w[153][47] = 5'b10000; w[153][48] = 5'b10000; w[153][49] = 5'b10000; w[153][50] = 5'b10000; w[153][51] = 5'b10000; w[153][52] = 5'b10000; w[153][53] = 5'b01111; w[153][54] = 5'b01111; w[153][55] = 5'b01111; w[153][56] = 5'b01111; w[153][57] = 5'b01111; w[153][58] = 5'b01111; w[153][59] = 5'b00000; w[153][60] = 5'b00000; w[153][61] = 5'b01111; w[153][62] = 5'b10000; w[153][63] = 5'b00000; w[153][64] = 5'b01111; w[153][65] = 5'b00000; w[153][66] = 5'b00000; w[153][67] = 5'b01111; w[153][68] = 5'b01111; w[153][69] = 5'b01111; w[153][70] = 5'b01111; w[153][71] = 5'b01111; w[153][72] = 5'b01111; w[153][73] = 5'b00000; w[153][74] = 5'b01111; w[153][75] = 5'b01111; w[153][76] = 5'b10000; w[153][77] = 5'b00000; w[153][78] = 5'b01111; w[153][79] = 5'b01111; w[153][80] = 5'b00000; w[153][81] = 5'b01111; w[153][82] = 5'b01111; w[153][83] = 5'b01111; w[153][84] = 5'b01111; w[153][85] = 5'b01111; w[153][86] = 5'b01111; w[153][87] = 5'b00000; w[153][88] = 5'b01111; w[153][89] = 5'b01111; w[153][90] = 5'b10000; w[153][91] = 5'b10000; w[153][92] = 5'b01111; w[153][93] = 5'b01111; w[153][94] = 5'b01111; w[153][95] = 5'b01111; w[153][96] = 5'b01111; w[153][97] = 5'b01111; w[153][98] = 5'b01111; w[153][99] = 5'b01111; w[153][100] = 5'b01111; w[153][101] = 5'b00000; w[153][102] = 5'b01111; w[153][103] = 5'b01111; w[153][104] = 5'b10000; w[153][105] = 5'b10000; w[153][106] = 5'b01111; w[153][107] = 5'b00000; w[153][108] = 5'b00000; w[153][109] = 5'b01111; w[153][110] = 5'b01111; w[153][111] = 5'b01111; w[153][112] = 5'b01111; w[153][113] = 5'b01111; w[153][114] = 5'b01111; w[153][115] = 5'b00000; w[153][116] = 5'b01111; w[153][117] = 5'b01111; w[153][118] = 5'b10000; w[153][119] = 5'b10000; w[153][120] = 5'b00000; w[153][121] = 5'b00000; w[153][122] = 5'b00000; w[153][123] = 5'b01111; w[153][124] = 5'b01111; w[153][125] = 5'b01111; w[153][126] = 5'b01111; w[153][127] = 5'b01111; w[153][128] = 5'b01111; w[153][129] = 5'b00000; w[153][130] = 5'b01111; w[153][131] = 5'b01111; w[153][132] = 5'b00000; w[153][133] = 5'b10000; w[153][134] = 5'b01111; w[153][135] = 5'b01111; w[153][136] = 5'b00000; w[153][137] = 5'b01111; w[153][138] = 5'b01111; w[153][139] = 5'b01111; w[153][140] = 5'b01111; w[153][141] = 5'b01111; w[153][142] = 5'b01111; w[153][143] = 5'b00000; w[153][144] = 5'b00000; w[153][145] = 5'b01111; w[153][146] = 5'b00000; w[153][147] = 5'b10000; w[153][148] = 5'b01111; w[153][149] = 5'b00000; w[153][150] = 5'b00000; w[153][151] = 5'b01111; w[153][152] = 5'b01111; w[153][153] = 5'b00000; w[153][154] = 5'b01111; w[153][155] = 5'b01111; w[153][156] = 5'b01111; w[153][157] = 5'b00000; w[153][158] = 5'b00000; w[153][159] = 5'b00000; w[153][160] = 5'b10000; w[153][161] = 5'b10000; w[153][162] = 5'b10000; w[153][163] = 5'b00000; w[153][164] = 5'b00000; w[153][165] = 5'b01111; w[153][166] = 5'b01111; w[153][167] = 5'b01111; w[153][168] = 5'b01111; w[153][169] = 5'b01111; w[153][170] = 5'b01111; w[153][171] = 5'b01111; w[153][172] = 5'b00000; w[153][173] = 5'b00000; w[153][174] = 5'b10000; w[153][175] = 5'b10000; w[153][176] = 5'b10000; w[153][177] = 5'b00000; w[153][178] = 5'b01111; w[153][179] = 5'b01111; w[153][180] = 5'b01111; w[153][181] = 5'b01111; w[153][182] = 5'b01111; w[153][183] = 5'b01111; w[153][184] = 5'b01111; w[153][185] = 5'b01111; w[153][186] = 5'b01111; w[153][187] = 5'b01111; w[153][188] = 5'b01111; w[153][189] = 5'b01111; w[153][190] = 5'b01111; w[153][191] = 5'b01111; w[153][192] = 5'b01111; w[153][193] = 5'b01111; w[153][194] = 5'b01111; w[153][195] = 5'b01111; w[153][196] = 5'b01111; w[153][197] = 5'b01111; w[153][198] = 5'b01111; w[153][199] = 5'b01111; w[153][200] = 5'b01111; w[153][201] = 5'b01111; w[153][202] = 5'b01111; w[153][203] = 5'b01111; w[153][204] = 5'b01111; w[153][205] = 5'b01111; w[153][206] = 5'b01111; w[153][207] = 5'b01111; w[153][208] = 5'b01111; w[153][209] = 5'b01111; 
w[154][0] = 5'b01111; w[154][1] = 5'b01111; w[154][2] = 5'b01111; w[154][3] = 5'b01111; w[154][4] = 5'b01111; w[154][5] = 5'b01111; w[154][6] = 5'b01111; w[154][7] = 5'b01111; w[154][8] = 5'b01111; w[154][9] = 5'b01111; w[154][10] = 5'b01111; w[154][11] = 5'b01111; w[154][12] = 5'b01111; w[154][13] = 5'b01111; w[154][14] = 5'b01111; w[154][15] = 5'b01111; w[154][16] = 5'b01111; w[154][17] = 5'b01111; w[154][18] = 5'b01111; w[154][19] = 5'b01111; w[154][20] = 5'b01111; w[154][21] = 5'b01111; w[154][22] = 5'b01111; w[154][23] = 5'b01111; w[154][24] = 5'b01111; w[154][25] = 5'b01111; w[154][26] = 5'b01111; w[154][27] = 5'b01111; w[154][28] = 5'b01111; w[154][29] = 5'b01111; w[154][30] = 5'b01111; w[154][31] = 5'b00000; w[154][32] = 5'b10000; w[154][33] = 5'b10000; w[154][34] = 5'b10000; w[154][35] = 5'b10000; w[154][36] = 5'b10000; w[154][37] = 5'b10000; w[154][38] = 5'b00000; w[154][39] = 5'b01111; w[154][40] = 5'b01111; w[154][41] = 5'b01111; w[154][42] = 5'b01111; w[154][43] = 5'b01111; w[154][44] = 5'b01111; w[154][45] = 5'b10000; w[154][46] = 5'b10000; w[154][47] = 5'b10000; w[154][48] = 5'b10000; w[154][49] = 5'b10000; w[154][50] = 5'b10000; w[154][51] = 5'b10000; w[154][52] = 5'b10000; w[154][53] = 5'b01111; w[154][54] = 5'b01111; w[154][55] = 5'b01111; w[154][56] = 5'b01111; w[154][57] = 5'b01111; w[154][58] = 5'b01111; w[154][59] = 5'b00000; w[154][60] = 5'b00000; w[154][61] = 5'b01111; w[154][62] = 5'b10000; w[154][63] = 5'b00000; w[154][64] = 5'b01111; w[154][65] = 5'b00000; w[154][66] = 5'b00000; w[154][67] = 5'b01111; w[154][68] = 5'b01111; w[154][69] = 5'b01111; w[154][70] = 5'b01111; w[154][71] = 5'b01111; w[154][72] = 5'b01111; w[154][73] = 5'b00000; w[154][74] = 5'b01111; w[154][75] = 5'b01111; w[154][76] = 5'b10000; w[154][77] = 5'b00000; w[154][78] = 5'b01111; w[154][79] = 5'b01111; w[154][80] = 5'b00000; w[154][81] = 5'b01111; w[154][82] = 5'b01111; w[154][83] = 5'b01111; w[154][84] = 5'b01111; w[154][85] = 5'b01111; w[154][86] = 5'b01111; w[154][87] = 5'b00000; w[154][88] = 5'b01111; w[154][89] = 5'b01111; w[154][90] = 5'b10000; w[154][91] = 5'b10000; w[154][92] = 5'b01111; w[154][93] = 5'b01111; w[154][94] = 5'b01111; w[154][95] = 5'b01111; w[154][96] = 5'b01111; w[154][97] = 5'b01111; w[154][98] = 5'b01111; w[154][99] = 5'b01111; w[154][100] = 5'b01111; w[154][101] = 5'b00000; w[154][102] = 5'b01111; w[154][103] = 5'b01111; w[154][104] = 5'b10000; w[154][105] = 5'b10000; w[154][106] = 5'b01111; w[154][107] = 5'b00000; w[154][108] = 5'b00000; w[154][109] = 5'b01111; w[154][110] = 5'b01111; w[154][111] = 5'b01111; w[154][112] = 5'b01111; w[154][113] = 5'b01111; w[154][114] = 5'b01111; w[154][115] = 5'b00000; w[154][116] = 5'b01111; w[154][117] = 5'b01111; w[154][118] = 5'b10000; w[154][119] = 5'b10000; w[154][120] = 5'b00000; w[154][121] = 5'b00000; w[154][122] = 5'b00000; w[154][123] = 5'b01111; w[154][124] = 5'b01111; w[154][125] = 5'b01111; w[154][126] = 5'b01111; w[154][127] = 5'b01111; w[154][128] = 5'b01111; w[154][129] = 5'b00000; w[154][130] = 5'b01111; w[154][131] = 5'b01111; w[154][132] = 5'b00000; w[154][133] = 5'b10000; w[154][134] = 5'b01111; w[154][135] = 5'b01111; w[154][136] = 5'b00000; w[154][137] = 5'b01111; w[154][138] = 5'b01111; w[154][139] = 5'b01111; w[154][140] = 5'b01111; w[154][141] = 5'b01111; w[154][142] = 5'b01111; w[154][143] = 5'b00000; w[154][144] = 5'b00000; w[154][145] = 5'b01111; w[154][146] = 5'b00000; w[154][147] = 5'b10000; w[154][148] = 5'b01111; w[154][149] = 5'b00000; w[154][150] = 5'b00000; w[154][151] = 5'b01111; w[154][152] = 5'b01111; w[154][153] = 5'b01111; w[154][154] = 5'b00000; w[154][155] = 5'b01111; w[154][156] = 5'b01111; w[154][157] = 5'b00000; w[154][158] = 5'b00000; w[154][159] = 5'b00000; w[154][160] = 5'b10000; w[154][161] = 5'b10000; w[154][162] = 5'b10000; w[154][163] = 5'b00000; w[154][164] = 5'b00000; w[154][165] = 5'b01111; w[154][166] = 5'b01111; w[154][167] = 5'b01111; w[154][168] = 5'b01111; w[154][169] = 5'b01111; w[154][170] = 5'b01111; w[154][171] = 5'b01111; w[154][172] = 5'b00000; w[154][173] = 5'b00000; w[154][174] = 5'b10000; w[154][175] = 5'b10000; w[154][176] = 5'b10000; w[154][177] = 5'b00000; w[154][178] = 5'b01111; w[154][179] = 5'b01111; w[154][180] = 5'b01111; w[154][181] = 5'b01111; w[154][182] = 5'b01111; w[154][183] = 5'b01111; w[154][184] = 5'b01111; w[154][185] = 5'b01111; w[154][186] = 5'b01111; w[154][187] = 5'b01111; w[154][188] = 5'b01111; w[154][189] = 5'b01111; w[154][190] = 5'b01111; w[154][191] = 5'b01111; w[154][192] = 5'b01111; w[154][193] = 5'b01111; w[154][194] = 5'b01111; w[154][195] = 5'b01111; w[154][196] = 5'b01111; w[154][197] = 5'b01111; w[154][198] = 5'b01111; w[154][199] = 5'b01111; w[154][200] = 5'b01111; w[154][201] = 5'b01111; w[154][202] = 5'b01111; w[154][203] = 5'b01111; w[154][204] = 5'b01111; w[154][205] = 5'b01111; w[154][206] = 5'b01111; w[154][207] = 5'b01111; w[154][208] = 5'b01111; w[154][209] = 5'b01111; 
w[155][0] = 5'b01111; w[155][1] = 5'b01111; w[155][2] = 5'b01111; w[155][3] = 5'b01111; w[155][4] = 5'b01111; w[155][5] = 5'b01111; w[155][6] = 5'b01111; w[155][7] = 5'b01111; w[155][8] = 5'b01111; w[155][9] = 5'b01111; w[155][10] = 5'b01111; w[155][11] = 5'b01111; w[155][12] = 5'b01111; w[155][13] = 5'b01111; w[155][14] = 5'b01111; w[155][15] = 5'b01111; w[155][16] = 5'b01111; w[155][17] = 5'b01111; w[155][18] = 5'b01111; w[155][19] = 5'b01111; w[155][20] = 5'b01111; w[155][21] = 5'b01111; w[155][22] = 5'b01111; w[155][23] = 5'b01111; w[155][24] = 5'b01111; w[155][25] = 5'b01111; w[155][26] = 5'b01111; w[155][27] = 5'b01111; w[155][28] = 5'b01111; w[155][29] = 5'b01111; w[155][30] = 5'b01111; w[155][31] = 5'b00000; w[155][32] = 5'b10000; w[155][33] = 5'b10000; w[155][34] = 5'b10000; w[155][35] = 5'b10000; w[155][36] = 5'b10000; w[155][37] = 5'b10000; w[155][38] = 5'b00000; w[155][39] = 5'b01111; w[155][40] = 5'b01111; w[155][41] = 5'b01111; w[155][42] = 5'b01111; w[155][43] = 5'b01111; w[155][44] = 5'b01111; w[155][45] = 5'b10000; w[155][46] = 5'b10000; w[155][47] = 5'b10000; w[155][48] = 5'b10000; w[155][49] = 5'b10000; w[155][50] = 5'b10000; w[155][51] = 5'b10000; w[155][52] = 5'b10000; w[155][53] = 5'b01111; w[155][54] = 5'b01111; w[155][55] = 5'b01111; w[155][56] = 5'b01111; w[155][57] = 5'b01111; w[155][58] = 5'b01111; w[155][59] = 5'b00000; w[155][60] = 5'b00000; w[155][61] = 5'b01111; w[155][62] = 5'b10000; w[155][63] = 5'b00000; w[155][64] = 5'b01111; w[155][65] = 5'b00000; w[155][66] = 5'b00000; w[155][67] = 5'b01111; w[155][68] = 5'b01111; w[155][69] = 5'b01111; w[155][70] = 5'b01111; w[155][71] = 5'b01111; w[155][72] = 5'b01111; w[155][73] = 5'b00000; w[155][74] = 5'b01111; w[155][75] = 5'b01111; w[155][76] = 5'b10000; w[155][77] = 5'b00000; w[155][78] = 5'b01111; w[155][79] = 5'b01111; w[155][80] = 5'b00000; w[155][81] = 5'b01111; w[155][82] = 5'b01111; w[155][83] = 5'b01111; w[155][84] = 5'b01111; w[155][85] = 5'b01111; w[155][86] = 5'b01111; w[155][87] = 5'b00000; w[155][88] = 5'b01111; w[155][89] = 5'b01111; w[155][90] = 5'b10000; w[155][91] = 5'b10000; w[155][92] = 5'b01111; w[155][93] = 5'b01111; w[155][94] = 5'b01111; w[155][95] = 5'b01111; w[155][96] = 5'b01111; w[155][97] = 5'b01111; w[155][98] = 5'b01111; w[155][99] = 5'b01111; w[155][100] = 5'b01111; w[155][101] = 5'b00000; w[155][102] = 5'b01111; w[155][103] = 5'b01111; w[155][104] = 5'b10000; w[155][105] = 5'b10000; w[155][106] = 5'b01111; w[155][107] = 5'b00000; w[155][108] = 5'b00000; w[155][109] = 5'b01111; w[155][110] = 5'b01111; w[155][111] = 5'b01111; w[155][112] = 5'b01111; w[155][113] = 5'b01111; w[155][114] = 5'b01111; w[155][115] = 5'b00000; w[155][116] = 5'b01111; w[155][117] = 5'b01111; w[155][118] = 5'b10000; w[155][119] = 5'b10000; w[155][120] = 5'b00000; w[155][121] = 5'b00000; w[155][122] = 5'b00000; w[155][123] = 5'b01111; w[155][124] = 5'b01111; w[155][125] = 5'b01111; w[155][126] = 5'b01111; w[155][127] = 5'b01111; w[155][128] = 5'b01111; w[155][129] = 5'b00000; w[155][130] = 5'b01111; w[155][131] = 5'b01111; w[155][132] = 5'b00000; w[155][133] = 5'b10000; w[155][134] = 5'b01111; w[155][135] = 5'b01111; w[155][136] = 5'b00000; w[155][137] = 5'b01111; w[155][138] = 5'b01111; w[155][139] = 5'b01111; w[155][140] = 5'b01111; w[155][141] = 5'b01111; w[155][142] = 5'b01111; w[155][143] = 5'b00000; w[155][144] = 5'b00000; w[155][145] = 5'b01111; w[155][146] = 5'b00000; w[155][147] = 5'b10000; w[155][148] = 5'b01111; w[155][149] = 5'b00000; w[155][150] = 5'b00000; w[155][151] = 5'b01111; w[155][152] = 5'b01111; w[155][153] = 5'b01111; w[155][154] = 5'b01111; w[155][155] = 5'b00000; w[155][156] = 5'b01111; w[155][157] = 5'b00000; w[155][158] = 5'b00000; w[155][159] = 5'b00000; w[155][160] = 5'b10000; w[155][161] = 5'b10000; w[155][162] = 5'b10000; w[155][163] = 5'b00000; w[155][164] = 5'b00000; w[155][165] = 5'b01111; w[155][166] = 5'b01111; w[155][167] = 5'b01111; w[155][168] = 5'b01111; w[155][169] = 5'b01111; w[155][170] = 5'b01111; w[155][171] = 5'b01111; w[155][172] = 5'b00000; w[155][173] = 5'b00000; w[155][174] = 5'b10000; w[155][175] = 5'b10000; w[155][176] = 5'b10000; w[155][177] = 5'b00000; w[155][178] = 5'b01111; w[155][179] = 5'b01111; w[155][180] = 5'b01111; w[155][181] = 5'b01111; w[155][182] = 5'b01111; w[155][183] = 5'b01111; w[155][184] = 5'b01111; w[155][185] = 5'b01111; w[155][186] = 5'b01111; w[155][187] = 5'b01111; w[155][188] = 5'b01111; w[155][189] = 5'b01111; w[155][190] = 5'b01111; w[155][191] = 5'b01111; w[155][192] = 5'b01111; w[155][193] = 5'b01111; w[155][194] = 5'b01111; w[155][195] = 5'b01111; w[155][196] = 5'b01111; w[155][197] = 5'b01111; w[155][198] = 5'b01111; w[155][199] = 5'b01111; w[155][200] = 5'b01111; w[155][201] = 5'b01111; w[155][202] = 5'b01111; w[155][203] = 5'b01111; w[155][204] = 5'b01111; w[155][205] = 5'b01111; w[155][206] = 5'b01111; w[155][207] = 5'b01111; w[155][208] = 5'b01111; w[155][209] = 5'b01111; 
w[156][0] = 5'b01111; w[156][1] = 5'b01111; w[156][2] = 5'b01111; w[156][3] = 5'b01111; w[156][4] = 5'b01111; w[156][5] = 5'b01111; w[156][6] = 5'b01111; w[156][7] = 5'b01111; w[156][8] = 5'b01111; w[156][9] = 5'b01111; w[156][10] = 5'b01111; w[156][11] = 5'b01111; w[156][12] = 5'b01111; w[156][13] = 5'b01111; w[156][14] = 5'b01111; w[156][15] = 5'b01111; w[156][16] = 5'b01111; w[156][17] = 5'b01111; w[156][18] = 5'b01111; w[156][19] = 5'b01111; w[156][20] = 5'b01111; w[156][21] = 5'b01111; w[156][22] = 5'b01111; w[156][23] = 5'b01111; w[156][24] = 5'b01111; w[156][25] = 5'b01111; w[156][26] = 5'b01111; w[156][27] = 5'b01111; w[156][28] = 5'b01111; w[156][29] = 5'b01111; w[156][30] = 5'b01111; w[156][31] = 5'b00000; w[156][32] = 5'b10000; w[156][33] = 5'b10000; w[156][34] = 5'b10000; w[156][35] = 5'b10000; w[156][36] = 5'b10000; w[156][37] = 5'b10000; w[156][38] = 5'b00000; w[156][39] = 5'b01111; w[156][40] = 5'b01111; w[156][41] = 5'b01111; w[156][42] = 5'b01111; w[156][43] = 5'b01111; w[156][44] = 5'b01111; w[156][45] = 5'b10000; w[156][46] = 5'b10000; w[156][47] = 5'b10000; w[156][48] = 5'b10000; w[156][49] = 5'b10000; w[156][50] = 5'b10000; w[156][51] = 5'b10000; w[156][52] = 5'b10000; w[156][53] = 5'b01111; w[156][54] = 5'b01111; w[156][55] = 5'b01111; w[156][56] = 5'b01111; w[156][57] = 5'b01111; w[156][58] = 5'b01111; w[156][59] = 5'b00000; w[156][60] = 5'b00000; w[156][61] = 5'b01111; w[156][62] = 5'b10000; w[156][63] = 5'b00000; w[156][64] = 5'b01111; w[156][65] = 5'b00000; w[156][66] = 5'b00000; w[156][67] = 5'b01111; w[156][68] = 5'b01111; w[156][69] = 5'b01111; w[156][70] = 5'b01111; w[156][71] = 5'b01111; w[156][72] = 5'b01111; w[156][73] = 5'b00000; w[156][74] = 5'b01111; w[156][75] = 5'b01111; w[156][76] = 5'b10000; w[156][77] = 5'b00000; w[156][78] = 5'b01111; w[156][79] = 5'b01111; w[156][80] = 5'b00000; w[156][81] = 5'b01111; w[156][82] = 5'b01111; w[156][83] = 5'b01111; w[156][84] = 5'b01111; w[156][85] = 5'b01111; w[156][86] = 5'b01111; w[156][87] = 5'b00000; w[156][88] = 5'b01111; w[156][89] = 5'b01111; w[156][90] = 5'b10000; w[156][91] = 5'b10000; w[156][92] = 5'b01111; w[156][93] = 5'b01111; w[156][94] = 5'b01111; w[156][95] = 5'b01111; w[156][96] = 5'b01111; w[156][97] = 5'b01111; w[156][98] = 5'b01111; w[156][99] = 5'b01111; w[156][100] = 5'b01111; w[156][101] = 5'b00000; w[156][102] = 5'b01111; w[156][103] = 5'b01111; w[156][104] = 5'b10000; w[156][105] = 5'b10000; w[156][106] = 5'b01111; w[156][107] = 5'b00000; w[156][108] = 5'b00000; w[156][109] = 5'b01111; w[156][110] = 5'b01111; w[156][111] = 5'b01111; w[156][112] = 5'b01111; w[156][113] = 5'b01111; w[156][114] = 5'b01111; w[156][115] = 5'b00000; w[156][116] = 5'b01111; w[156][117] = 5'b01111; w[156][118] = 5'b10000; w[156][119] = 5'b10000; w[156][120] = 5'b00000; w[156][121] = 5'b00000; w[156][122] = 5'b00000; w[156][123] = 5'b01111; w[156][124] = 5'b01111; w[156][125] = 5'b01111; w[156][126] = 5'b01111; w[156][127] = 5'b01111; w[156][128] = 5'b01111; w[156][129] = 5'b00000; w[156][130] = 5'b01111; w[156][131] = 5'b01111; w[156][132] = 5'b00000; w[156][133] = 5'b10000; w[156][134] = 5'b01111; w[156][135] = 5'b01111; w[156][136] = 5'b00000; w[156][137] = 5'b01111; w[156][138] = 5'b01111; w[156][139] = 5'b01111; w[156][140] = 5'b01111; w[156][141] = 5'b01111; w[156][142] = 5'b01111; w[156][143] = 5'b00000; w[156][144] = 5'b00000; w[156][145] = 5'b01111; w[156][146] = 5'b00000; w[156][147] = 5'b10000; w[156][148] = 5'b01111; w[156][149] = 5'b00000; w[156][150] = 5'b00000; w[156][151] = 5'b01111; w[156][152] = 5'b01111; w[156][153] = 5'b01111; w[156][154] = 5'b01111; w[156][155] = 5'b01111; w[156][156] = 5'b00000; w[156][157] = 5'b00000; w[156][158] = 5'b00000; w[156][159] = 5'b00000; w[156][160] = 5'b10000; w[156][161] = 5'b10000; w[156][162] = 5'b10000; w[156][163] = 5'b00000; w[156][164] = 5'b00000; w[156][165] = 5'b01111; w[156][166] = 5'b01111; w[156][167] = 5'b01111; w[156][168] = 5'b01111; w[156][169] = 5'b01111; w[156][170] = 5'b01111; w[156][171] = 5'b01111; w[156][172] = 5'b00000; w[156][173] = 5'b00000; w[156][174] = 5'b10000; w[156][175] = 5'b10000; w[156][176] = 5'b10000; w[156][177] = 5'b00000; w[156][178] = 5'b01111; w[156][179] = 5'b01111; w[156][180] = 5'b01111; w[156][181] = 5'b01111; w[156][182] = 5'b01111; w[156][183] = 5'b01111; w[156][184] = 5'b01111; w[156][185] = 5'b01111; w[156][186] = 5'b01111; w[156][187] = 5'b01111; w[156][188] = 5'b01111; w[156][189] = 5'b01111; w[156][190] = 5'b01111; w[156][191] = 5'b01111; w[156][192] = 5'b01111; w[156][193] = 5'b01111; w[156][194] = 5'b01111; w[156][195] = 5'b01111; w[156][196] = 5'b01111; w[156][197] = 5'b01111; w[156][198] = 5'b01111; w[156][199] = 5'b01111; w[156][200] = 5'b01111; w[156][201] = 5'b01111; w[156][202] = 5'b01111; w[156][203] = 5'b01111; w[156][204] = 5'b01111; w[156][205] = 5'b01111; w[156][206] = 5'b01111; w[156][207] = 5'b01111; w[156][208] = 5'b01111; w[156][209] = 5'b01111; 
w[157][0] = 5'b00000; w[157][1] = 5'b00000; w[157][2] = 5'b00000; w[157][3] = 5'b00000; w[157][4] = 5'b00000; w[157][5] = 5'b00000; w[157][6] = 5'b00000; w[157][7] = 5'b00000; w[157][8] = 5'b00000; w[157][9] = 5'b00000; w[157][10] = 5'b00000; w[157][11] = 5'b00000; w[157][12] = 5'b00000; w[157][13] = 5'b00000; w[157][14] = 5'b00000; w[157][15] = 5'b00000; w[157][16] = 5'b00000; w[157][17] = 5'b00000; w[157][18] = 5'b00000; w[157][19] = 5'b00000; w[157][20] = 5'b00000; w[157][21] = 5'b00000; w[157][22] = 5'b00000; w[157][23] = 5'b00000; w[157][24] = 5'b00000; w[157][25] = 5'b00000; w[157][26] = 5'b00000; w[157][27] = 5'b00000; w[157][28] = 5'b00000; w[157][29] = 5'b00000; w[157][30] = 5'b10000; w[157][31] = 5'b00000; w[157][32] = 5'b01111; w[157][33] = 5'b00000; w[157][34] = 5'b10000; w[157][35] = 5'b10000; w[157][36] = 5'b10000; w[157][37] = 5'b01111; w[157][38] = 5'b00000; w[157][39] = 5'b10000; w[157][40] = 5'b00000; w[157][41] = 5'b00000; w[157][42] = 5'b00000; w[157][43] = 5'b00000; w[157][44] = 5'b10000; w[157][45] = 5'b01111; w[157][46] = 5'b01111; w[157][47] = 5'b00000; w[157][48] = 5'b10000; w[157][49] = 5'b10000; w[157][50] = 5'b10000; w[157][51] = 5'b01111; w[157][52] = 5'b01111; w[157][53] = 5'b10000; w[157][54] = 5'b00000; w[157][55] = 5'b00000; w[157][56] = 5'b00000; w[157][57] = 5'b00000; w[157][58] = 5'b01111; w[157][59] = 5'b01111; w[157][60] = 5'b01111; w[157][61] = 5'b01111; w[157][62] = 5'b10000; w[157][63] = 5'b10000; w[157][64] = 5'b00000; w[157][65] = 5'b01111; w[157][66] = 5'b01111; w[157][67] = 5'b01111; w[157][68] = 5'b00000; w[157][69] = 5'b00000; w[157][70] = 5'b00000; w[157][71] = 5'b00000; w[157][72] = 5'b01111; w[157][73] = 5'b01111; w[157][74] = 5'b01111; w[157][75] = 5'b01111; w[157][76] = 5'b10000; w[157][77] = 5'b10000; w[157][78] = 5'b00000; w[157][79] = 5'b01111; w[157][80] = 5'b01111; w[157][81] = 5'b01111; w[157][82] = 5'b00000; w[157][83] = 5'b00000; w[157][84] = 5'b00000; w[157][85] = 5'b00000; w[157][86] = 5'b01111; w[157][87] = 5'b01111; w[157][88] = 5'b01111; w[157][89] = 5'b01111; w[157][90] = 5'b10000; w[157][91] = 5'b10000; w[157][92] = 5'b00000; w[157][93] = 5'b01111; w[157][94] = 5'b01111; w[157][95] = 5'b00000; w[157][96] = 5'b00000; w[157][97] = 5'b00000; w[157][98] = 5'b00000; w[157][99] = 5'b00000; w[157][100] = 5'b01111; w[157][101] = 5'b01111; w[157][102] = 5'b01111; w[157][103] = 5'b00000; w[157][104] = 5'b10000; w[157][105] = 5'b10000; w[157][106] = 5'b01111; w[157][107] = 5'b01111; w[157][108] = 5'b01111; w[157][109] = 5'b01111; w[157][110] = 5'b00000; w[157][111] = 5'b00000; w[157][112] = 5'b00000; w[157][113] = 5'b00000; w[157][114] = 5'b01111; w[157][115] = 5'b01111; w[157][116] = 5'b01111; w[157][117] = 5'b00000; w[157][118] = 5'b10000; w[157][119] = 5'b10000; w[157][120] = 5'b01111; w[157][121] = 5'b01111; w[157][122] = 5'b01111; w[157][123] = 5'b01111; w[157][124] = 5'b00000; w[157][125] = 5'b00000; w[157][126] = 5'b00000; w[157][127] = 5'b00000; w[157][128] = 5'b01111; w[157][129] = 5'b01111; w[157][130] = 5'b01111; w[157][131] = 5'b00000; w[157][132] = 5'b10000; w[157][133] = 5'b10000; w[157][134] = 5'b01111; w[157][135] = 5'b01111; w[157][136] = 5'b01111; w[157][137] = 5'b01111; w[157][138] = 5'b00000; w[157][139] = 5'b00000; w[157][140] = 5'b00000; w[157][141] = 5'b00000; w[157][142] = 5'b01111; w[157][143] = 5'b01111; w[157][144] = 5'b01111; w[157][145] = 5'b00000; w[157][146] = 5'b10000; w[157][147] = 5'b10000; w[157][148] = 5'b01111; w[157][149] = 5'b01111; w[157][150] = 5'b01111; w[157][151] = 5'b01111; w[157][152] = 5'b00000; w[157][153] = 5'b00000; w[157][154] = 5'b00000; w[157][155] = 5'b00000; w[157][156] = 5'b00000; w[157][157] = 5'b00000; w[157][158] = 5'b01111; w[157][159] = 5'b00000; w[157][160] = 5'b10000; w[157][161] = 5'b10000; w[157][162] = 5'b01111; w[157][163] = 5'b01111; w[157][164] = 5'b01111; w[157][165] = 5'b00000; w[157][166] = 5'b00000; w[157][167] = 5'b00000; w[157][168] = 5'b00000; w[157][169] = 5'b00000; w[157][170] = 5'b00000; w[157][171] = 5'b01111; w[157][172] = 5'b01111; w[157][173] = 5'b00000; w[157][174] = 5'b10000; w[157][175] = 5'b10000; w[157][176] = 5'b01111; w[157][177] = 5'b01111; w[157][178] = 5'b01111; w[157][179] = 5'b00000; w[157][180] = 5'b00000; w[157][181] = 5'b00000; w[157][182] = 5'b00000; w[157][183] = 5'b00000; w[157][184] = 5'b00000; w[157][185] = 5'b00000; w[157][186] = 5'b00000; w[157][187] = 5'b00000; w[157][188] = 5'b00000; w[157][189] = 5'b00000; w[157][190] = 5'b00000; w[157][191] = 5'b00000; w[157][192] = 5'b00000; w[157][193] = 5'b00000; w[157][194] = 5'b00000; w[157][195] = 5'b00000; w[157][196] = 5'b00000; w[157][197] = 5'b00000; w[157][198] = 5'b00000; w[157][199] = 5'b00000; w[157][200] = 5'b00000; w[157][201] = 5'b00000; w[157][202] = 5'b00000; w[157][203] = 5'b00000; w[157][204] = 5'b00000; w[157][205] = 5'b00000; w[157][206] = 5'b00000; w[157][207] = 5'b00000; w[157][208] = 5'b00000; w[157][209] = 5'b00000; 
w[158][0] = 5'b00000; w[158][1] = 5'b00000; w[158][2] = 5'b00000; w[158][3] = 5'b00000; w[158][4] = 5'b00000; w[158][5] = 5'b00000; w[158][6] = 5'b00000; w[158][7] = 5'b00000; w[158][8] = 5'b00000; w[158][9] = 5'b00000; w[158][10] = 5'b00000; w[158][11] = 5'b00000; w[158][12] = 5'b00000; w[158][13] = 5'b00000; w[158][14] = 5'b00000; w[158][15] = 5'b00000; w[158][16] = 5'b00000; w[158][17] = 5'b00000; w[158][18] = 5'b00000; w[158][19] = 5'b00000; w[158][20] = 5'b00000; w[158][21] = 5'b00000; w[158][22] = 5'b00000; w[158][23] = 5'b00000; w[158][24] = 5'b00000; w[158][25] = 5'b00000; w[158][26] = 5'b00000; w[158][27] = 5'b00000; w[158][28] = 5'b00000; w[158][29] = 5'b00000; w[158][30] = 5'b10000; w[158][31] = 5'b00000; w[158][32] = 5'b01111; w[158][33] = 5'b00000; w[158][34] = 5'b10000; w[158][35] = 5'b10000; w[158][36] = 5'b10000; w[158][37] = 5'b01111; w[158][38] = 5'b00000; w[158][39] = 5'b10000; w[158][40] = 5'b00000; w[158][41] = 5'b00000; w[158][42] = 5'b00000; w[158][43] = 5'b00000; w[158][44] = 5'b10000; w[158][45] = 5'b01111; w[158][46] = 5'b01111; w[158][47] = 5'b00000; w[158][48] = 5'b10000; w[158][49] = 5'b10000; w[158][50] = 5'b10000; w[158][51] = 5'b01111; w[158][52] = 5'b01111; w[158][53] = 5'b10000; w[158][54] = 5'b00000; w[158][55] = 5'b00000; w[158][56] = 5'b00000; w[158][57] = 5'b00000; w[158][58] = 5'b01111; w[158][59] = 5'b01111; w[158][60] = 5'b01111; w[158][61] = 5'b01111; w[158][62] = 5'b10000; w[158][63] = 5'b10000; w[158][64] = 5'b00000; w[158][65] = 5'b01111; w[158][66] = 5'b01111; w[158][67] = 5'b01111; w[158][68] = 5'b00000; w[158][69] = 5'b00000; w[158][70] = 5'b00000; w[158][71] = 5'b00000; w[158][72] = 5'b01111; w[158][73] = 5'b01111; w[158][74] = 5'b01111; w[158][75] = 5'b01111; w[158][76] = 5'b10000; w[158][77] = 5'b10000; w[158][78] = 5'b00000; w[158][79] = 5'b01111; w[158][80] = 5'b01111; w[158][81] = 5'b01111; w[158][82] = 5'b00000; w[158][83] = 5'b00000; w[158][84] = 5'b00000; w[158][85] = 5'b00000; w[158][86] = 5'b01111; w[158][87] = 5'b01111; w[158][88] = 5'b01111; w[158][89] = 5'b01111; w[158][90] = 5'b10000; w[158][91] = 5'b10000; w[158][92] = 5'b00000; w[158][93] = 5'b01111; w[158][94] = 5'b01111; w[158][95] = 5'b00000; w[158][96] = 5'b00000; w[158][97] = 5'b00000; w[158][98] = 5'b00000; w[158][99] = 5'b00000; w[158][100] = 5'b01111; w[158][101] = 5'b01111; w[158][102] = 5'b01111; w[158][103] = 5'b00000; w[158][104] = 5'b10000; w[158][105] = 5'b10000; w[158][106] = 5'b01111; w[158][107] = 5'b01111; w[158][108] = 5'b01111; w[158][109] = 5'b01111; w[158][110] = 5'b00000; w[158][111] = 5'b00000; w[158][112] = 5'b00000; w[158][113] = 5'b00000; w[158][114] = 5'b01111; w[158][115] = 5'b01111; w[158][116] = 5'b01111; w[158][117] = 5'b00000; w[158][118] = 5'b10000; w[158][119] = 5'b10000; w[158][120] = 5'b01111; w[158][121] = 5'b01111; w[158][122] = 5'b01111; w[158][123] = 5'b01111; w[158][124] = 5'b00000; w[158][125] = 5'b00000; w[158][126] = 5'b00000; w[158][127] = 5'b00000; w[158][128] = 5'b01111; w[158][129] = 5'b01111; w[158][130] = 5'b01111; w[158][131] = 5'b00000; w[158][132] = 5'b10000; w[158][133] = 5'b10000; w[158][134] = 5'b01111; w[158][135] = 5'b01111; w[158][136] = 5'b01111; w[158][137] = 5'b01111; w[158][138] = 5'b00000; w[158][139] = 5'b00000; w[158][140] = 5'b00000; w[158][141] = 5'b00000; w[158][142] = 5'b01111; w[158][143] = 5'b01111; w[158][144] = 5'b01111; w[158][145] = 5'b00000; w[158][146] = 5'b10000; w[158][147] = 5'b10000; w[158][148] = 5'b01111; w[158][149] = 5'b01111; w[158][150] = 5'b01111; w[158][151] = 5'b01111; w[158][152] = 5'b00000; w[158][153] = 5'b00000; w[158][154] = 5'b00000; w[158][155] = 5'b00000; w[158][156] = 5'b00000; w[158][157] = 5'b01111; w[158][158] = 5'b00000; w[158][159] = 5'b00000; w[158][160] = 5'b10000; w[158][161] = 5'b10000; w[158][162] = 5'b01111; w[158][163] = 5'b01111; w[158][164] = 5'b01111; w[158][165] = 5'b00000; w[158][166] = 5'b00000; w[158][167] = 5'b00000; w[158][168] = 5'b00000; w[158][169] = 5'b00000; w[158][170] = 5'b00000; w[158][171] = 5'b01111; w[158][172] = 5'b01111; w[158][173] = 5'b00000; w[158][174] = 5'b10000; w[158][175] = 5'b10000; w[158][176] = 5'b01111; w[158][177] = 5'b01111; w[158][178] = 5'b01111; w[158][179] = 5'b00000; w[158][180] = 5'b00000; w[158][181] = 5'b00000; w[158][182] = 5'b00000; w[158][183] = 5'b00000; w[158][184] = 5'b00000; w[158][185] = 5'b00000; w[158][186] = 5'b00000; w[158][187] = 5'b00000; w[158][188] = 5'b00000; w[158][189] = 5'b00000; w[158][190] = 5'b00000; w[158][191] = 5'b00000; w[158][192] = 5'b00000; w[158][193] = 5'b00000; w[158][194] = 5'b00000; w[158][195] = 5'b00000; w[158][196] = 5'b00000; w[158][197] = 5'b00000; w[158][198] = 5'b00000; w[158][199] = 5'b00000; w[158][200] = 5'b00000; w[158][201] = 5'b00000; w[158][202] = 5'b00000; w[158][203] = 5'b00000; w[158][204] = 5'b00000; w[158][205] = 5'b00000; w[158][206] = 5'b00000; w[158][207] = 5'b00000; w[158][208] = 5'b00000; w[158][209] = 5'b00000; 
w[159][0] = 5'b00000; w[159][1] = 5'b00000; w[159][2] = 5'b00000; w[159][3] = 5'b00000; w[159][4] = 5'b00000; w[159][5] = 5'b00000; w[159][6] = 5'b00000; w[159][7] = 5'b00000; w[159][8] = 5'b00000; w[159][9] = 5'b00000; w[159][10] = 5'b00000; w[159][11] = 5'b00000; w[159][12] = 5'b00000; w[159][13] = 5'b00000; w[159][14] = 5'b00000; w[159][15] = 5'b00000; w[159][16] = 5'b00000; w[159][17] = 5'b00000; w[159][18] = 5'b00000; w[159][19] = 5'b00000; w[159][20] = 5'b00000; w[159][21] = 5'b00000; w[159][22] = 5'b00000; w[159][23] = 5'b00000; w[159][24] = 5'b00000; w[159][25] = 5'b00000; w[159][26] = 5'b00000; w[159][27] = 5'b00000; w[159][28] = 5'b00000; w[159][29] = 5'b00000; w[159][30] = 5'b10000; w[159][31] = 5'b10000; w[159][32] = 5'b10000; w[159][33] = 5'b00000; w[159][34] = 5'b01111; w[159][35] = 5'b01111; w[159][36] = 5'b01111; w[159][37] = 5'b10000; w[159][38] = 5'b10000; w[159][39] = 5'b10000; w[159][40] = 5'b00000; w[159][41] = 5'b00000; w[159][42] = 5'b00000; w[159][43] = 5'b00000; w[159][44] = 5'b10000; w[159][45] = 5'b10000; w[159][46] = 5'b10000; w[159][47] = 5'b00000; w[159][48] = 5'b01111; w[159][49] = 5'b01111; w[159][50] = 5'b01111; w[159][51] = 5'b10000; w[159][52] = 5'b10000; w[159][53] = 5'b10000; w[159][54] = 5'b00000; w[159][55] = 5'b00000; w[159][56] = 5'b00000; w[159][57] = 5'b00000; w[159][58] = 5'b01111; w[159][59] = 5'b00000; w[159][60] = 5'b00000; w[159][61] = 5'b10000; w[159][62] = 5'b10000; w[159][63] = 5'b00000; w[159][64] = 5'b00000; w[159][65] = 5'b00000; w[159][66] = 5'b00000; w[159][67] = 5'b01111; w[159][68] = 5'b00000; w[159][69] = 5'b00000; w[159][70] = 5'b00000; w[159][71] = 5'b00000; w[159][72] = 5'b01111; w[159][73] = 5'b00000; w[159][74] = 5'b10000; w[159][75] = 5'b10000; w[159][76] = 5'b10000; w[159][77] = 5'b00000; w[159][78] = 5'b00000; w[159][79] = 5'b10000; w[159][80] = 5'b00000; w[159][81] = 5'b01111; w[159][82] = 5'b00000; w[159][83] = 5'b00000; w[159][84] = 5'b00000; w[159][85] = 5'b00000; w[159][86] = 5'b01111; w[159][87] = 5'b00000; w[159][88] = 5'b10000; w[159][89] = 5'b10000; w[159][90] = 5'b10000; w[159][91] = 5'b10000; w[159][92] = 5'b00000; w[159][93] = 5'b10000; w[159][94] = 5'b10000; w[159][95] = 5'b00000; w[159][96] = 5'b00000; w[159][97] = 5'b00000; w[159][98] = 5'b00000; w[159][99] = 5'b00000; w[159][100] = 5'b01111; w[159][101] = 5'b00000; w[159][102] = 5'b10000; w[159][103] = 5'b00000; w[159][104] = 5'b10000; w[159][105] = 5'b10000; w[159][106] = 5'b01111; w[159][107] = 5'b00000; w[159][108] = 5'b00000; w[159][109] = 5'b01111; w[159][110] = 5'b00000; w[159][111] = 5'b00000; w[159][112] = 5'b00000; w[159][113] = 5'b00000; w[159][114] = 5'b01111; w[159][115] = 5'b00000; w[159][116] = 5'b10000; w[159][117] = 5'b00000; w[159][118] = 5'b10000; w[159][119] = 5'b10000; w[159][120] = 5'b00000; w[159][121] = 5'b00000; w[159][122] = 5'b00000; w[159][123] = 5'b01111; w[159][124] = 5'b00000; w[159][125] = 5'b00000; w[159][126] = 5'b00000; w[159][127] = 5'b00000; w[159][128] = 5'b01111; w[159][129] = 5'b00000; w[159][130] = 5'b10000; w[159][131] = 5'b00000; w[159][132] = 5'b00000; w[159][133] = 5'b10000; w[159][134] = 5'b10000; w[159][135] = 5'b10000; w[159][136] = 5'b00000; w[159][137] = 5'b01111; w[159][138] = 5'b00000; w[159][139] = 5'b00000; w[159][140] = 5'b00000; w[159][141] = 5'b00000; w[159][142] = 5'b01111; w[159][143] = 5'b00000; w[159][144] = 5'b00000; w[159][145] = 5'b00000; w[159][146] = 5'b00000; w[159][147] = 5'b10000; w[159][148] = 5'b10000; w[159][149] = 5'b00000; w[159][150] = 5'b00000; w[159][151] = 5'b01111; w[159][152] = 5'b00000; w[159][153] = 5'b00000; w[159][154] = 5'b00000; w[159][155] = 5'b00000; w[159][156] = 5'b00000; w[159][157] = 5'b00000; w[159][158] = 5'b00000; w[159][159] = 5'b00000; w[159][160] = 5'b01111; w[159][161] = 5'b01111; w[159][162] = 5'b01111; w[159][163] = 5'b00000; w[159][164] = 5'b00000; w[159][165] = 5'b00000; w[159][166] = 5'b00000; w[159][167] = 5'b00000; w[159][168] = 5'b00000; w[159][169] = 5'b00000; w[159][170] = 5'b00000; w[159][171] = 5'b10000; w[159][172] = 5'b00000; w[159][173] = 5'b01111; w[159][174] = 5'b01111; w[159][175] = 5'b01111; w[159][176] = 5'b01111; w[159][177] = 5'b00000; w[159][178] = 5'b10000; w[159][179] = 5'b00000; w[159][180] = 5'b00000; w[159][181] = 5'b00000; w[159][182] = 5'b00000; w[159][183] = 5'b00000; w[159][184] = 5'b00000; w[159][185] = 5'b00000; w[159][186] = 5'b00000; w[159][187] = 5'b00000; w[159][188] = 5'b00000; w[159][189] = 5'b00000; w[159][190] = 5'b00000; w[159][191] = 5'b00000; w[159][192] = 5'b00000; w[159][193] = 5'b00000; w[159][194] = 5'b00000; w[159][195] = 5'b00000; w[159][196] = 5'b00000; w[159][197] = 5'b00000; w[159][198] = 5'b00000; w[159][199] = 5'b00000; w[159][200] = 5'b00000; w[159][201] = 5'b00000; w[159][202] = 5'b00000; w[159][203] = 5'b00000; w[159][204] = 5'b00000; w[159][205] = 5'b00000; w[159][206] = 5'b00000; w[159][207] = 5'b00000; w[159][208] = 5'b00000; w[159][209] = 5'b00000; 
w[160][0] = 5'b10000; w[160][1] = 5'b10000; w[160][2] = 5'b10000; w[160][3] = 5'b10000; w[160][4] = 5'b10000; w[160][5] = 5'b10000; w[160][6] = 5'b10000; w[160][7] = 5'b10000; w[160][8] = 5'b10000; w[160][9] = 5'b10000; w[160][10] = 5'b10000; w[160][11] = 5'b10000; w[160][12] = 5'b10000; w[160][13] = 5'b10000; w[160][14] = 5'b10000; w[160][15] = 5'b10000; w[160][16] = 5'b10000; w[160][17] = 5'b10000; w[160][18] = 5'b10000; w[160][19] = 5'b10000; w[160][20] = 5'b10000; w[160][21] = 5'b10000; w[160][22] = 5'b10000; w[160][23] = 5'b10000; w[160][24] = 5'b10000; w[160][25] = 5'b10000; w[160][26] = 5'b10000; w[160][27] = 5'b10000; w[160][28] = 5'b10000; w[160][29] = 5'b10000; w[160][30] = 5'b00000; w[160][31] = 5'b10000; w[160][32] = 5'b00000; w[160][33] = 5'b01111; w[160][34] = 5'b01111; w[160][35] = 5'b01111; w[160][36] = 5'b01111; w[160][37] = 5'b00000; w[160][38] = 5'b10000; w[160][39] = 5'b00000; w[160][40] = 5'b10000; w[160][41] = 5'b10000; w[160][42] = 5'b10000; w[160][43] = 5'b10000; w[160][44] = 5'b00000; w[160][45] = 5'b00000; w[160][46] = 5'b00000; w[160][47] = 5'b01111; w[160][48] = 5'b01111; w[160][49] = 5'b01111; w[160][50] = 5'b01111; w[160][51] = 5'b00000; w[160][52] = 5'b00000; w[160][53] = 5'b00000; w[160][54] = 5'b10000; w[160][55] = 5'b10000; w[160][56] = 5'b10000; w[160][57] = 5'b10000; w[160][58] = 5'b00000; w[160][59] = 5'b10000; w[160][60] = 5'b10000; w[160][61] = 5'b10000; w[160][62] = 5'b00000; w[160][63] = 5'b01111; w[160][64] = 5'b10000; w[160][65] = 5'b10000; w[160][66] = 5'b10000; w[160][67] = 5'b00000; w[160][68] = 5'b10000; w[160][69] = 5'b10000; w[160][70] = 5'b10000; w[160][71] = 5'b10000; w[160][72] = 5'b00000; w[160][73] = 5'b10000; w[160][74] = 5'b10000; w[160][75] = 5'b10000; w[160][76] = 5'b00000; w[160][77] = 5'b01111; w[160][78] = 5'b10000; w[160][79] = 5'b10000; w[160][80] = 5'b10000; w[160][81] = 5'b00000; w[160][82] = 5'b10000; w[160][83] = 5'b10000; w[160][84] = 5'b10000; w[160][85] = 5'b10000; w[160][86] = 5'b00000; w[160][87] = 5'b10000; w[160][88] = 5'b10000; w[160][89] = 5'b10000; w[160][90] = 5'b00000; w[160][91] = 5'b00000; w[160][92] = 5'b10000; w[160][93] = 5'b10000; w[160][94] = 5'b10000; w[160][95] = 5'b10000; w[160][96] = 5'b10000; w[160][97] = 5'b10000; w[160][98] = 5'b10000; w[160][99] = 5'b10000; w[160][100] = 5'b00000; w[160][101] = 5'b10000; w[160][102] = 5'b10000; w[160][103] = 5'b10000; w[160][104] = 5'b00000; w[160][105] = 5'b00000; w[160][106] = 5'b00000; w[160][107] = 5'b10000; w[160][108] = 5'b10000; w[160][109] = 5'b00000; w[160][110] = 5'b10000; w[160][111] = 5'b10000; w[160][112] = 5'b10000; w[160][113] = 5'b10000; w[160][114] = 5'b00000; w[160][115] = 5'b10000; w[160][116] = 5'b10000; w[160][117] = 5'b10000; w[160][118] = 5'b00000; w[160][119] = 5'b00000; w[160][120] = 5'b10000; w[160][121] = 5'b10000; w[160][122] = 5'b10000; w[160][123] = 5'b00000; w[160][124] = 5'b10000; w[160][125] = 5'b10000; w[160][126] = 5'b10000; w[160][127] = 5'b10000; w[160][128] = 5'b00000; w[160][129] = 5'b10000; w[160][130] = 5'b10000; w[160][131] = 5'b10000; w[160][132] = 5'b01111; w[160][133] = 5'b00000; w[160][134] = 5'b10000; w[160][135] = 5'b10000; w[160][136] = 5'b10000; w[160][137] = 5'b00000; w[160][138] = 5'b10000; w[160][139] = 5'b10000; w[160][140] = 5'b10000; w[160][141] = 5'b10000; w[160][142] = 5'b00000; w[160][143] = 5'b10000; w[160][144] = 5'b10000; w[160][145] = 5'b10000; w[160][146] = 5'b01111; w[160][147] = 5'b00000; w[160][148] = 5'b10000; w[160][149] = 5'b10000; w[160][150] = 5'b10000; w[160][151] = 5'b00000; w[160][152] = 5'b10000; w[160][153] = 5'b10000; w[160][154] = 5'b10000; w[160][155] = 5'b10000; w[160][156] = 5'b10000; w[160][157] = 5'b10000; w[160][158] = 5'b10000; w[160][159] = 5'b01111; w[160][160] = 5'b00000; w[160][161] = 5'b01111; w[160][162] = 5'b00000; w[160][163] = 5'b10000; w[160][164] = 5'b10000; w[160][165] = 5'b10000; w[160][166] = 5'b10000; w[160][167] = 5'b10000; w[160][168] = 5'b10000; w[160][169] = 5'b10000; w[160][170] = 5'b10000; w[160][171] = 5'b10000; w[160][172] = 5'b10000; w[160][173] = 5'b01111; w[160][174] = 5'b01111; w[160][175] = 5'b01111; w[160][176] = 5'b00000; w[160][177] = 5'b10000; w[160][178] = 5'b10000; w[160][179] = 5'b10000; w[160][180] = 5'b10000; w[160][181] = 5'b10000; w[160][182] = 5'b10000; w[160][183] = 5'b10000; w[160][184] = 5'b10000; w[160][185] = 5'b10000; w[160][186] = 5'b10000; w[160][187] = 5'b10000; w[160][188] = 5'b10000; w[160][189] = 5'b10000; w[160][190] = 5'b10000; w[160][191] = 5'b10000; w[160][192] = 5'b10000; w[160][193] = 5'b10000; w[160][194] = 5'b10000; w[160][195] = 5'b10000; w[160][196] = 5'b10000; w[160][197] = 5'b10000; w[160][198] = 5'b10000; w[160][199] = 5'b10000; w[160][200] = 5'b10000; w[160][201] = 5'b10000; w[160][202] = 5'b10000; w[160][203] = 5'b10000; w[160][204] = 5'b10000; w[160][205] = 5'b10000; w[160][206] = 5'b10000; w[160][207] = 5'b10000; w[160][208] = 5'b10000; w[160][209] = 5'b10000; 
w[161][0] = 5'b10000; w[161][1] = 5'b10000; w[161][2] = 5'b10000; w[161][3] = 5'b10000; w[161][4] = 5'b10000; w[161][5] = 5'b10000; w[161][6] = 5'b10000; w[161][7] = 5'b10000; w[161][8] = 5'b10000; w[161][9] = 5'b10000; w[161][10] = 5'b10000; w[161][11] = 5'b10000; w[161][12] = 5'b10000; w[161][13] = 5'b10000; w[161][14] = 5'b10000; w[161][15] = 5'b10000; w[161][16] = 5'b10000; w[161][17] = 5'b10000; w[161][18] = 5'b10000; w[161][19] = 5'b10000; w[161][20] = 5'b10000; w[161][21] = 5'b10000; w[161][22] = 5'b10000; w[161][23] = 5'b10000; w[161][24] = 5'b10000; w[161][25] = 5'b10000; w[161][26] = 5'b10000; w[161][27] = 5'b10000; w[161][28] = 5'b10000; w[161][29] = 5'b10000; w[161][30] = 5'b00000; w[161][31] = 5'b10000; w[161][32] = 5'b00000; w[161][33] = 5'b01111; w[161][34] = 5'b01111; w[161][35] = 5'b01111; w[161][36] = 5'b01111; w[161][37] = 5'b00000; w[161][38] = 5'b10000; w[161][39] = 5'b00000; w[161][40] = 5'b10000; w[161][41] = 5'b10000; w[161][42] = 5'b10000; w[161][43] = 5'b10000; w[161][44] = 5'b00000; w[161][45] = 5'b00000; w[161][46] = 5'b00000; w[161][47] = 5'b01111; w[161][48] = 5'b01111; w[161][49] = 5'b01111; w[161][50] = 5'b01111; w[161][51] = 5'b00000; w[161][52] = 5'b00000; w[161][53] = 5'b00000; w[161][54] = 5'b10000; w[161][55] = 5'b10000; w[161][56] = 5'b10000; w[161][57] = 5'b10000; w[161][58] = 5'b00000; w[161][59] = 5'b10000; w[161][60] = 5'b10000; w[161][61] = 5'b10000; w[161][62] = 5'b00000; w[161][63] = 5'b01111; w[161][64] = 5'b10000; w[161][65] = 5'b10000; w[161][66] = 5'b10000; w[161][67] = 5'b00000; w[161][68] = 5'b10000; w[161][69] = 5'b10000; w[161][70] = 5'b10000; w[161][71] = 5'b10000; w[161][72] = 5'b00000; w[161][73] = 5'b10000; w[161][74] = 5'b10000; w[161][75] = 5'b10000; w[161][76] = 5'b00000; w[161][77] = 5'b01111; w[161][78] = 5'b10000; w[161][79] = 5'b10000; w[161][80] = 5'b10000; w[161][81] = 5'b00000; w[161][82] = 5'b10000; w[161][83] = 5'b10000; w[161][84] = 5'b10000; w[161][85] = 5'b10000; w[161][86] = 5'b00000; w[161][87] = 5'b10000; w[161][88] = 5'b10000; w[161][89] = 5'b10000; w[161][90] = 5'b00000; w[161][91] = 5'b00000; w[161][92] = 5'b10000; w[161][93] = 5'b10000; w[161][94] = 5'b10000; w[161][95] = 5'b10000; w[161][96] = 5'b10000; w[161][97] = 5'b10000; w[161][98] = 5'b10000; w[161][99] = 5'b10000; w[161][100] = 5'b00000; w[161][101] = 5'b10000; w[161][102] = 5'b10000; w[161][103] = 5'b10000; w[161][104] = 5'b00000; w[161][105] = 5'b00000; w[161][106] = 5'b00000; w[161][107] = 5'b10000; w[161][108] = 5'b10000; w[161][109] = 5'b00000; w[161][110] = 5'b10000; w[161][111] = 5'b10000; w[161][112] = 5'b10000; w[161][113] = 5'b10000; w[161][114] = 5'b00000; w[161][115] = 5'b10000; w[161][116] = 5'b10000; w[161][117] = 5'b10000; w[161][118] = 5'b00000; w[161][119] = 5'b00000; w[161][120] = 5'b10000; w[161][121] = 5'b10000; w[161][122] = 5'b10000; w[161][123] = 5'b00000; w[161][124] = 5'b10000; w[161][125] = 5'b10000; w[161][126] = 5'b10000; w[161][127] = 5'b10000; w[161][128] = 5'b00000; w[161][129] = 5'b10000; w[161][130] = 5'b10000; w[161][131] = 5'b10000; w[161][132] = 5'b01111; w[161][133] = 5'b00000; w[161][134] = 5'b10000; w[161][135] = 5'b10000; w[161][136] = 5'b10000; w[161][137] = 5'b00000; w[161][138] = 5'b10000; w[161][139] = 5'b10000; w[161][140] = 5'b10000; w[161][141] = 5'b10000; w[161][142] = 5'b00000; w[161][143] = 5'b10000; w[161][144] = 5'b10000; w[161][145] = 5'b10000; w[161][146] = 5'b01111; w[161][147] = 5'b00000; w[161][148] = 5'b10000; w[161][149] = 5'b10000; w[161][150] = 5'b10000; w[161][151] = 5'b00000; w[161][152] = 5'b10000; w[161][153] = 5'b10000; w[161][154] = 5'b10000; w[161][155] = 5'b10000; w[161][156] = 5'b10000; w[161][157] = 5'b10000; w[161][158] = 5'b10000; w[161][159] = 5'b01111; w[161][160] = 5'b01111; w[161][161] = 5'b00000; w[161][162] = 5'b00000; w[161][163] = 5'b10000; w[161][164] = 5'b10000; w[161][165] = 5'b10000; w[161][166] = 5'b10000; w[161][167] = 5'b10000; w[161][168] = 5'b10000; w[161][169] = 5'b10000; w[161][170] = 5'b10000; w[161][171] = 5'b10000; w[161][172] = 5'b10000; w[161][173] = 5'b01111; w[161][174] = 5'b01111; w[161][175] = 5'b01111; w[161][176] = 5'b00000; w[161][177] = 5'b10000; w[161][178] = 5'b10000; w[161][179] = 5'b10000; w[161][180] = 5'b10000; w[161][181] = 5'b10000; w[161][182] = 5'b10000; w[161][183] = 5'b10000; w[161][184] = 5'b10000; w[161][185] = 5'b10000; w[161][186] = 5'b10000; w[161][187] = 5'b10000; w[161][188] = 5'b10000; w[161][189] = 5'b10000; w[161][190] = 5'b10000; w[161][191] = 5'b10000; w[161][192] = 5'b10000; w[161][193] = 5'b10000; w[161][194] = 5'b10000; w[161][195] = 5'b10000; w[161][196] = 5'b10000; w[161][197] = 5'b10000; w[161][198] = 5'b10000; w[161][199] = 5'b10000; w[161][200] = 5'b10000; w[161][201] = 5'b10000; w[161][202] = 5'b10000; w[161][203] = 5'b10000; w[161][204] = 5'b10000; w[161][205] = 5'b10000; w[161][206] = 5'b10000; w[161][207] = 5'b10000; w[161][208] = 5'b10000; w[161][209] = 5'b10000; 
w[162][0] = 5'b10000; w[162][1] = 5'b10000; w[162][2] = 5'b10000; w[162][3] = 5'b10000; w[162][4] = 5'b10000; w[162][5] = 5'b10000; w[162][6] = 5'b10000; w[162][7] = 5'b10000; w[162][8] = 5'b10000; w[162][9] = 5'b10000; w[162][10] = 5'b10000; w[162][11] = 5'b10000; w[162][12] = 5'b10000; w[162][13] = 5'b10000; w[162][14] = 5'b10000; w[162][15] = 5'b10000; w[162][16] = 5'b10000; w[162][17] = 5'b10000; w[162][18] = 5'b10000; w[162][19] = 5'b10000; w[162][20] = 5'b10000; w[162][21] = 5'b10000; w[162][22] = 5'b10000; w[162][23] = 5'b10000; w[162][24] = 5'b10000; w[162][25] = 5'b10000; w[162][26] = 5'b10000; w[162][27] = 5'b10000; w[162][28] = 5'b10000; w[162][29] = 5'b10000; w[162][30] = 5'b10000; w[162][31] = 5'b10000; w[162][32] = 5'b00000; w[162][33] = 5'b01111; w[162][34] = 5'b00000; w[162][35] = 5'b00000; w[162][36] = 5'b00000; w[162][37] = 5'b00000; w[162][38] = 5'b10000; w[162][39] = 5'b10000; w[162][40] = 5'b10000; w[162][41] = 5'b10000; w[162][42] = 5'b10000; w[162][43] = 5'b10000; w[162][44] = 5'b10000; w[162][45] = 5'b00000; w[162][46] = 5'b00000; w[162][47] = 5'b01111; w[162][48] = 5'b00000; w[162][49] = 5'b00000; w[162][50] = 5'b00000; w[162][51] = 5'b00000; w[162][52] = 5'b00000; w[162][53] = 5'b10000; w[162][54] = 5'b10000; w[162][55] = 5'b10000; w[162][56] = 5'b10000; w[162][57] = 5'b10000; w[162][58] = 5'b00000; w[162][59] = 5'b01111; w[162][60] = 5'b01111; w[162][61] = 5'b00000; w[162][62] = 5'b00000; w[162][63] = 5'b10000; w[162][64] = 5'b10000; w[162][65] = 5'b01111; w[162][66] = 5'b01111; w[162][67] = 5'b00000; w[162][68] = 5'b10000; w[162][69] = 5'b10000; w[162][70] = 5'b10000; w[162][71] = 5'b10000; w[162][72] = 5'b00000; w[162][73] = 5'b01111; w[162][74] = 5'b00000; w[162][75] = 5'b00000; w[162][76] = 5'b00000; w[162][77] = 5'b10000; w[162][78] = 5'b10000; w[162][79] = 5'b00000; w[162][80] = 5'b01111; w[162][81] = 5'b00000; w[162][82] = 5'b10000; w[162][83] = 5'b10000; w[162][84] = 5'b10000; w[162][85] = 5'b10000; w[162][86] = 5'b00000; w[162][87] = 5'b01111; w[162][88] = 5'b00000; w[162][89] = 5'b00000; w[162][90] = 5'b00000; w[162][91] = 5'b00000; w[162][92] = 5'b10000; w[162][93] = 5'b00000; w[162][94] = 5'b00000; w[162][95] = 5'b10000; w[162][96] = 5'b10000; w[162][97] = 5'b10000; w[162][98] = 5'b10000; w[162][99] = 5'b10000; w[162][100] = 5'b00000; w[162][101] = 5'b01111; w[162][102] = 5'b00000; w[162][103] = 5'b10000; w[162][104] = 5'b00000; w[162][105] = 5'b00000; w[162][106] = 5'b00000; w[162][107] = 5'b01111; w[162][108] = 5'b01111; w[162][109] = 5'b00000; w[162][110] = 5'b10000; w[162][111] = 5'b10000; w[162][112] = 5'b10000; w[162][113] = 5'b10000; w[162][114] = 5'b00000; w[162][115] = 5'b01111; w[162][116] = 5'b00000; w[162][117] = 5'b10000; w[162][118] = 5'b00000; w[162][119] = 5'b00000; w[162][120] = 5'b01111; w[162][121] = 5'b01111; w[162][122] = 5'b01111; w[162][123] = 5'b00000; w[162][124] = 5'b10000; w[162][125] = 5'b10000; w[162][126] = 5'b10000; w[162][127] = 5'b10000; w[162][128] = 5'b00000; w[162][129] = 5'b01111; w[162][130] = 5'b00000; w[162][131] = 5'b10000; w[162][132] = 5'b10000; w[162][133] = 5'b00000; w[162][134] = 5'b00000; w[162][135] = 5'b00000; w[162][136] = 5'b01111; w[162][137] = 5'b00000; w[162][138] = 5'b10000; w[162][139] = 5'b10000; w[162][140] = 5'b10000; w[162][141] = 5'b10000; w[162][142] = 5'b00000; w[162][143] = 5'b01111; w[162][144] = 5'b01111; w[162][145] = 5'b10000; w[162][146] = 5'b10000; w[162][147] = 5'b00000; w[162][148] = 5'b00000; w[162][149] = 5'b01111; w[162][150] = 5'b01111; w[162][151] = 5'b00000; w[162][152] = 5'b10000; w[162][153] = 5'b10000; w[162][154] = 5'b10000; w[162][155] = 5'b10000; w[162][156] = 5'b10000; w[162][157] = 5'b01111; w[162][158] = 5'b01111; w[162][159] = 5'b01111; w[162][160] = 5'b00000; w[162][161] = 5'b00000; w[162][162] = 5'b00000; w[162][163] = 5'b01111; w[162][164] = 5'b01111; w[162][165] = 5'b10000; w[162][166] = 5'b10000; w[162][167] = 5'b10000; w[162][168] = 5'b10000; w[162][169] = 5'b10000; w[162][170] = 5'b10000; w[162][171] = 5'b00000; w[162][172] = 5'b01111; w[162][173] = 5'b01111; w[162][174] = 5'b00000; w[162][175] = 5'b00000; w[162][176] = 5'b01111; w[162][177] = 5'b01111; w[162][178] = 5'b00000; w[162][179] = 5'b10000; w[162][180] = 5'b10000; w[162][181] = 5'b10000; w[162][182] = 5'b10000; w[162][183] = 5'b10000; w[162][184] = 5'b10000; w[162][185] = 5'b10000; w[162][186] = 5'b10000; w[162][187] = 5'b10000; w[162][188] = 5'b10000; w[162][189] = 5'b10000; w[162][190] = 5'b10000; w[162][191] = 5'b10000; w[162][192] = 5'b10000; w[162][193] = 5'b10000; w[162][194] = 5'b10000; w[162][195] = 5'b10000; w[162][196] = 5'b10000; w[162][197] = 5'b10000; w[162][198] = 5'b10000; w[162][199] = 5'b10000; w[162][200] = 5'b10000; w[162][201] = 5'b10000; w[162][202] = 5'b10000; w[162][203] = 5'b10000; w[162][204] = 5'b10000; w[162][205] = 5'b10000; w[162][206] = 5'b10000; w[162][207] = 5'b10000; w[162][208] = 5'b10000; w[162][209] = 5'b10000; 
w[163][0] = 5'b00000; w[163][1] = 5'b00000; w[163][2] = 5'b00000; w[163][3] = 5'b00000; w[163][4] = 5'b00000; w[163][5] = 5'b00000; w[163][6] = 5'b00000; w[163][7] = 5'b00000; w[163][8] = 5'b00000; w[163][9] = 5'b00000; w[163][10] = 5'b00000; w[163][11] = 5'b00000; w[163][12] = 5'b00000; w[163][13] = 5'b00000; w[163][14] = 5'b00000; w[163][15] = 5'b00000; w[163][16] = 5'b00000; w[163][17] = 5'b00000; w[163][18] = 5'b00000; w[163][19] = 5'b00000; w[163][20] = 5'b00000; w[163][21] = 5'b00000; w[163][22] = 5'b00000; w[163][23] = 5'b00000; w[163][24] = 5'b00000; w[163][25] = 5'b00000; w[163][26] = 5'b00000; w[163][27] = 5'b00000; w[163][28] = 5'b00000; w[163][29] = 5'b00000; w[163][30] = 5'b10000; w[163][31] = 5'b00000; w[163][32] = 5'b01111; w[163][33] = 5'b00000; w[163][34] = 5'b10000; w[163][35] = 5'b10000; w[163][36] = 5'b10000; w[163][37] = 5'b01111; w[163][38] = 5'b00000; w[163][39] = 5'b10000; w[163][40] = 5'b00000; w[163][41] = 5'b00000; w[163][42] = 5'b00000; w[163][43] = 5'b00000; w[163][44] = 5'b10000; w[163][45] = 5'b01111; w[163][46] = 5'b01111; w[163][47] = 5'b00000; w[163][48] = 5'b10000; w[163][49] = 5'b10000; w[163][50] = 5'b10000; w[163][51] = 5'b01111; w[163][52] = 5'b01111; w[163][53] = 5'b10000; w[163][54] = 5'b00000; w[163][55] = 5'b00000; w[163][56] = 5'b00000; w[163][57] = 5'b00000; w[163][58] = 5'b01111; w[163][59] = 5'b01111; w[163][60] = 5'b01111; w[163][61] = 5'b01111; w[163][62] = 5'b10000; w[163][63] = 5'b10000; w[163][64] = 5'b00000; w[163][65] = 5'b01111; w[163][66] = 5'b01111; w[163][67] = 5'b01111; w[163][68] = 5'b00000; w[163][69] = 5'b00000; w[163][70] = 5'b00000; w[163][71] = 5'b00000; w[163][72] = 5'b01111; w[163][73] = 5'b01111; w[163][74] = 5'b01111; w[163][75] = 5'b01111; w[163][76] = 5'b10000; w[163][77] = 5'b10000; w[163][78] = 5'b00000; w[163][79] = 5'b01111; w[163][80] = 5'b01111; w[163][81] = 5'b01111; w[163][82] = 5'b00000; w[163][83] = 5'b00000; w[163][84] = 5'b00000; w[163][85] = 5'b00000; w[163][86] = 5'b01111; w[163][87] = 5'b01111; w[163][88] = 5'b01111; w[163][89] = 5'b01111; w[163][90] = 5'b10000; w[163][91] = 5'b10000; w[163][92] = 5'b00000; w[163][93] = 5'b01111; w[163][94] = 5'b01111; w[163][95] = 5'b00000; w[163][96] = 5'b00000; w[163][97] = 5'b00000; w[163][98] = 5'b00000; w[163][99] = 5'b00000; w[163][100] = 5'b01111; w[163][101] = 5'b01111; w[163][102] = 5'b01111; w[163][103] = 5'b00000; w[163][104] = 5'b10000; w[163][105] = 5'b10000; w[163][106] = 5'b01111; w[163][107] = 5'b01111; w[163][108] = 5'b01111; w[163][109] = 5'b01111; w[163][110] = 5'b00000; w[163][111] = 5'b00000; w[163][112] = 5'b00000; w[163][113] = 5'b00000; w[163][114] = 5'b01111; w[163][115] = 5'b01111; w[163][116] = 5'b01111; w[163][117] = 5'b00000; w[163][118] = 5'b10000; w[163][119] = 5'b10000; w[163][120] = 5'b01111; w[163][121] = 5'b01111; w[163][122] = 5'b01111; w[163][123] = 5'b01111; w[163][124] = 5'b00000; w[163][125] = 5'b00000; w[163][126] = 5'b00000; w[163][127] = 5'b00000; w[163][128] = 5'b01111; w[163][129] = 5'b01111; w[163][130] = 5'b01111; w[163][131] = 5'b00000; w[163][132] = 5'b10000; w[163][133] = 5'b10000; w[163][134] = 5'b01111; w[163][135] = 5'b01111; w[163][136] = 5'b01111; w[163][137] = 5'b01111; w[163][138] = 5'b00000; w[163][139] = 5'b00000; w[163][140] = 5'b00000; w[163][141] = 5'b00000; w[163][142] = 5'b01111; w[163][143] = 5'b01111; w[163][144] = 5'b01111; w[163][145] = 5'b00000; w[163][146] = 5'b10000; w[163][147] = 5'b10000; w[163][148] = 5'b01111; w[163][149] = 5'b01111; w[163][150] = 5'b01111; w[163][151] = 5'b01111; w[163][152] = 5'b00000; w[163][153] = 5'b00000; w[163][154] = 5'b00000; w[163][155] = 5'b00000; w[163][156] = 5'b00000; w[163][157] = 5'b01111; w[163][158] = 5'b01111; w[163][159] = 5'b00000; w[163][160] = 5'b10000; w[163][161] = 5'b10000; w[163][162] = 5'b01111; w[163][163] = 5'b00000; w[163][164] = 5'b01111; w[163][165] = 5'b00000; w[163][166] = 5'b00000; w[163][167] = 5'b00000; w[163][168] = 5'b00000; w[163][169] = 5'b00000; w[163][170] = 5'b00000; w[163][171] = 5'b01111; w[163][172] = 5'b01111; w[163][173] = 5'b00000; w[163][174] = 5'b10000; w[163][175] = 5'b10000; w[163][176] = 5'b01111; w[163][177] = 5'b01111; w[163][178] = 5'b01111; w[163][179] = 5'b00000; w[163][180] = 5'b00000; w[163][181] = 5'b00000; w[163][182] = 5'b00000; w[163][183] = 5'b00000; w[163][184] = 5'b00000; w[163][185] = 5'b00000; w[163][186] = 5'b00000; w[163][187] = 5'b00000; w[163][188] = 5'b00000; w[163][189] = 5'b00000; w[163][190] = 5'b00000; w[163][191] = 5'b00000; w[163][192] = 5'b00000; w[163][193] = 5'b00000; w[163][194] = 5'b00000; w[163][195] = 5'b00000; w[163][196] = 5'b00000; w[163][197] = 5'b00000; w[163][198] = 5'b00000; w[163][199] = 5'b00000; w[163][200] = 5'b00000; w[163][201] = 5'b00000; w[163][202] = 5'b00000; w[163][203] = 5'b00000; w[163][204] = 5'b00000; w[163][205] = 5'b00000; w[163][206] = 5'b00000; w[163][207] = 5'b00000; w[163][208] = 5'b00000; w[163][209] = 5'b00000; 
w[164][0] = 5'b00000; w[164][1] = 5'b00000; w[164][2] = 5'b00000; w[164][3] = 5'b00000; w[164][4] = 5'b00000; w[164][5] = 5'b00000; w[164][6] = 5'b00000; w[164][7] = 5'b00000; w[164][8] = 5'b00000; w[164][9] = 5'b00000; w[164][10] = 5'b00000; w[164][11] = 5'b00000; w[164][12] = 5'b00000; w[164][13] = 5'b00000; w[164][14] = 5'b00000; w[164][15] = 5'b00000; w[164][16] = 5'b00000; w[164][17] = 5'b00000; w[164][18] = 5'b00000; w[164][19] = 5'b00000; w[164][20] = 5'b00000; w[164][21] = 5'b00000; w[164][22] = 5'b00000; w[164][23] = 5'b00000; w[164][24] = 5'b00000; w[164][25] = 5'b00000; w[164][26] = 5'b00000; w[164][27] = 5'b00000; w[164][28] = 5'b00000; w[164][29] = 5'b00000; w[164][30] = 5'b10000; w[164][31] = 5'b00000; w[164][32] = 5'b01111; w[164][33] = 5'b00000; w[164][34] = 5'b10000; w[164][35] = 5'b10000; w[164][36] = 5'b10000; w[164][37] = 5'b01111; w[164][38] = 5'b00000; w[164][39] = 5'b10000; w[164][40] = 5'b00000; w[164][41] = 5'b00000; w[164][42] = 5'b00000; w[164][43] = 5'b00000; w[164][44] = 5'b10000; w[164][45] = 5'b01111; w[164][46] = 5'b01111; w[164][47] = 5'b00000; w[164][48] = 5'b10000; w[164][49] = 5'b10000; w[164][50] = 5'b10000; w[164][51] = 5'b01111; w[164][52] = 5'b01111; w[164][53] = 5'b10000; w[164][54] = 5'b00000; w[164][55] = 5'b00000; w[164][56] = 5'b00000; w[164][57] = 5'b00000; w[164][58] = 5'b01111; w[164][59] = 5'b01111; w[164][60] = 5'b01111; w[164][61] = 5'b01111; w[164][62] = 5'b10000; w[164][63] = 5'b10000; w[164][64] = 5'b00000; w[164][65] = 5'b01111; w[164][66] = 5'b01111; w[164][67] = 5'b01111; w[164][68] = 5'b00000; w[164][69] = 5'b00000; w[164][70] = 5'b00000; w[164][71] = 5'b00000; w[164][72] = 5'b01111; w[164][73] = 5'b01111; w[164][74] = 5'b01111; w[164][75] = 5'b01111; w[164][76] = 5'b10000; w[164][77] = 5'b10000; w[164][78] = 5'b00000; w[164][79] = 5'b01111; w[164][80] = 5'b01111; w[164][81] = 5'b01111; w[164][82] = 5'b00000; w[164][83] = 5'b00000; w[164][84] = 5'b00000; w[164][85] = 5'b00000; w[164][86] = 5'b01111; w[164][87] = 5'b01111; w[164][88] = 5'b01111; w[164][89] = 5'b01111; w[164][90] = 5'b10000; w[164][91] = 5'b10000; w[164][92] = 5'b00000; w[164][93] = 5'b01111; w[164][94] = 5'b01111; w[164][95] = 5'b00000; w[164][96] = 5'b00000; w[164][97] = 5'b00000; w[164][98] = 5'b00000; w[164][99] = 5'b00000; w[164][100] = 5'b01111; w[164][101] = 5'b01111; w[164][102] = 5'b01111; w[164][103] = 5'b00000; w[164][104] = 5'b10000; w[164][105] = 5'b10000; w[164][106] = 5'b01111; w[164][107] = 5'b01111; w[164][108] = 5'b01111; w[164][109] = 5'b01111; w[164][110] = 5'b00000; w[164][111] = 5'b00000; w[164][112] = 5'b00000; w[164][113] = 5'b00000; w[164][114] = 5'b01111; w[164][115] = 5'b01111; w[164][116] = 5'b01111; w[164][117] = 5'b00000; w[164][118] = 5'b10000; w[164][119] = 5'b10000; w[164][120] = 5'b01111; w[164][121] = 5'b01111; w[164][122] = 5'b01111; w[164][123] = 5'b01111; w[164][124] = 5'b00000; w[164][125] = 5'b00000; w[164][126] = 5'b00000; w[164][127] = 5'b00000; w[164][128] = 5'b01111; w[164][129] = 5'b01111; w[164][130] = 5'b01111; w[164][131] = 5'b00000; w[164][132] = 5'b10000; w[164][133] = 5'b10000; w[164][134] = 5'b01111; w[164][135] = 5'b01111; w[164][136] = 5'b01111; w[164][137] = 5'b01111; w[164][138] = 5'b00000; w[164][139] = 5'b00000; w[164][140] = 5'b00000; w[164][141] = 5'b00000; w[164][142] = 5'b01111; w[164][143] = 5'b01111; w[164][144] = 5'b01111; w[164][145] = 5'b00000; w[164][146] = 5'b10000; w[164][147] = 5'b10000; w[164][148] = 5'b01111; w[164][149] = 5'b01111; w[164][150] = 5'b01111; w[164][151] = 5'b01111; w[164][152] = 5'b00000; w[164][153] = 5'b00000; w[164][154] = 5'b00000; w[164][155] = 5'b00000; w[164][156] = 5'b00000; w[164][157] = 5'b01111; w[164][158] = 5'b01111; w[164][159] = 5'b00000; w[164][160] = 5'b10000; w[164][161] = 5'b10000; w[164][162] = 5'b01111; w[164][163] = 5'b01111; w[164][164] = 5'b00000; w[164][165] = 5'b00000; w[164][166] = 5'b00000; w[164][167] = 5'b00000; w[164][168] = 5'b00000; w[164][169] = 5'b00000; w[164][170] = 5'b00000; w[164][171] = 5'b01111; w[164][172] = 5'b01111; w[164][173] = 5'b00000; w[164][174] = 5'b10000; w[164][175] = 5'b10000; w[164][176] = 5'b01111; w[164][177] = 5'b01111; w[164][178] = 5'b01111; w[164][179] = 5'b00000; w[164][180] = 5'b00000; w[164][181] = 5'b00000; w[164][182] = 5'b00000; w[164][183] = 5'b00000; w[164][184] = 5'b00000; w[164][185] = 5'b00000; w[164][186] = 5'b00000; w[164][187] = 5'b00000; w[164][188] = 5'b00000; w[164][189] = 5'b00000; w[164][190] = 5'b00000; w[164][191] = 5'b00000; w[164][192] = 5'b00000; w[164][193] = 5'b00000; w[164][194] = 5'b00000; w[164][195] = 5'b00000; w[164][196] = 5'b00000; w[164][197] = 5'b00000; w[164][198] = 5'b00000; w[164][199] = 5'b00000; w[164][200] = 5'b00000; w[164][201] = 5'b00000; w[164][202] = 5'b00000; w[164][203] = 5'b00000; w[164][204] = 5'b00000; w[164][205] = 5'b00000; w[164][206] = 5'b00000; w[164][207] = 5'b00000; w[164][208] = 5'b00000; w[164][209] = 5'b00000; 
w[165][0] = 5'b01111; w[165][1] = 5'b01111; w[165][2] = 5'b01111; w[165][3] = 5'b01111; w[165][4] = 5'b01111; w[165][5] = 5'b01111; w[165][6] = 5'b01111; w[165][7] = 5'b01111; w[165][8] = 5'b01111; w[165][9] = 5'b01111; w[165][10] = 5'b01111; w[165][11] = 5'b01111; w[165][12] = 5'b01111; w[165][13] = 5'b01111; w[165][14] = 5'b01111; w[165][15] = 5'b01111; w[165][16] = 5'b01111; w[165][17] = 5'b01111; w[165][18] = 5'b01111; w[165][19] = 5'b01111; w[165][20] = 5'b01111; w[165][21] = 5'b01111; w[165][22] = 5'b01111; w[165][23] = 5'b01111; w[165][24] = 5'b01111; w[165][25] = 5'b01111; w[165][26] = 5'b01111; w[165][27] = 5'b01111; w[165][28] = 5'b01111; w[165][29] = 5'b01111; w[165][30] = 5'b01111; w[165][31] = 5'b00000; w[165][32] = 5'b10000; w[165][33] = 5'b10000; w[165][34] = 5'b10000; w[165][35] = 5'b10000; w[165][36] = 5'b10000; w[165][37] = 5'b10000; w[165][38] = 5'b00000; w[165][39] = 5'b01111; w[165][40] = 5'b01111; w[165][41] = 5'b01111; w[165][42] = 5'b01111; w[165][43] = 5'b01111; w[165][44] = 5'b01111; w[165][45] = 5'b10000; w[165][46] = 5'b10000; w[165][47] = 5'b10000; w[165][48] = 5'b10000; w[165][49] = 5'b10000; w[165][50] = 5'b10000; w[165][51] = 5'b10000; w[165][52] = 5'b10000; w[165][53] = 5'b01111; w[165][54] = 5'b01111; w[165][55] = 5'b01111; w[165][56] = 5'b01111; w[165][57] = 5'b01111; w[165][58] = 5'b01111; w[165][59] = 5'b00000; w[165][60] = 5'b00000; w[165][61] = 5'b01111; w[165][62] = 5'b10000; w[165][63] = 5'b00000; w[165][64] = 5'b01111; w[165][65] = 5'b00000; w[165][66] = 5'b00000; w[165][67] = 5'b01111; w[165][68] = 5'b01111; w[165][69] = 5'b01111; w[165][70] = 5'b01111; w[165][71] = 5'b01111; w[165][72] = 5'b01111; w[165][73] = 5'b00000; w[165][74] = 5'b01111; w[165][75] = 5'b01111; w[165][76] = 5'b10000; w[165][77] = 5'b00000; w[165][78] = 5'b01111; w[165][79] = 5'b01111; w[165][80] = 5'b00000; w[165][81] = 5'b01111; w[165][82] = 5'b01111; w[165][83] = 5'b01111; w[165][84] = 5'b01111; w[165][85] = 5'b01111; w[165][86] = 5'b01111; w[165][87] = 5'b00000; w[165][88] = 5'b01111; w[165][89] = 5'b01111; w[165][90] = 5'b10000; w[165][91] = 5'b10000; w[165][92] = 5'b01111; w[165][93] = 5'b01111; w[165][94] = 5'b01111; w[165][95] = 5'b01111; w[165][96] = 5'b01111; w[165][97] = 5'b01111; w[165][98] = 5'b01111; w[165][99] = 5'b01111; w[165][100] = 5'b01111; w[165][101] = 5'b00000; w[165][102] = 5'b01111; w[165][103] = 5'b01111; w[165][104] = 5'b10000; w[165][105] = 5'b10000; w[165][106] = 5'b01111; w[165][107] = 5'b00000; w[165][108] = 5'b00000; w[165][109] = 5'b01111; w[165][110] = 5'b01111; w[165][111] = 5'b01111; w[165][112] = 5'b01111; w[165][113] = 5'b01111; w[165][114] = 5'b01111; w[165][115] = 5'b00000; w[165][116] = 5'b01111; w[165][117] = 5'b01111; w[165][118] = 5'b10000; w[165][119] = 5'b10000; w[165][120] = 5'b00000; w[165][121] = 5'b00000; w[165][122] = 5'b00000; w[165][123] = 5'b01111; w[165][124] = 5'b01111; w[165][125] = 5'b01111; w[165][126] = 5'b01111; w[165][127] = 5'b01111; w[165][128] = 5'b01111; w[165][129] = 5'b00000; w[165][130] = 5'b01111; w[165][131] = 5'b01111; w[165][132] = 5'b00000; w[165][133] = 5'b10000; w[165][134] = 5'b01111; w[165][135] = 5'b01111; w[165][136] = 5'b00000; w[165][137] = 5'b01111; w[165][138] = 5'b01111; w[165][139] = 5'b01111; w[165][140] = 5'b01111; w[165][141] = 5'b01111; w[165][142] = 5'b01111; w[165][143] = 5'b00000; w[165][144] = 5'b00000; w[165][145] = 5'b01111; w[165][146] = 5'b00000; w[165][147] = 5'b10000; w[165][148] = 5'b01111; w[165][149] = 5'b00000; w[165][150] = 5'b00000; w[165][151] = 5'b01111; w[165][152] = 5'b01111; w[165][153] = 5'b01111; w[165][154] = 5'b01111; w[165][155] = 5'b01111; w[165][156] = 5'b01111; w[165][157] = 5'b00000; w[165][158] = 5'b00000; w[165][159] = 5'b00000; w[165][160] = 5'b10000; w[165][161] = 5'b10000; w[165][162] = 5'b10000; w[165][163] = 5'b00000; w[165][164] = 5'b00000; w[165][165] = 5'b00000; w[165][166] = 5'b01111; w[165][167] = 5'b01111; w[165][168] = 5'b01111; w[165][169] = 5'b01111; w[165][170] = 5'b01111; w[165][171] = 5'b01111; w[165][172] = 5'b00000; w[165][173] = 5'b00000; w[165][174] = 5'b10000; w[165][175] = 5'b10000; w[165][176] = 5'b10000; w[165][177] = 5'b00000; w[165][178] = 5'b01111; w[165][179] = 5'b01111; w[165][180] = 5'b01111; w[165][181] = 5'b01111; w[165][182] = 5'b01111; w[165][183] = 5'b01111; w[165][184] = 5'b01111; w[165][185] = 5'b01111; w[165][186] = 5'b01111; w[165][187] = 5'b01111; w[165][188] = 5'b01111; w[165][189] = 5'b01111; w[165][190] = 5'b01111; w[165][191] = 5'b01111; w[165][192] = 5'b01111; w[165][193] = 5'b01111; w[165][194] = 5'b01111; w[165][195] = 5'b01111; w[165][196] = 5'b01111; w[165][197] = 5'b01111; w[165][198] = 5'b01111; w[165][199] = 5'b01111; w[165][200] = 5'b01111; w[165][201] = 5'b01111; w[165][202] = 5'b01111; w[165][203] = 5'b01111; w[165][204] = 5'b01111; w[165][205] = 5'b01111; w[165][206] = 5'b01111; w[165][207] = 5'b01111; w[165][208] = 5'b01111; w[165][209] = 5'b01111; 
w[166][0] = 5'b01111; w[166][1] = 5'b01111; w[166][2] = 5'b01111; w[166][3] = 5'b01111; w[166][4] = 5'b01111; w[166][5] = 5'b01111; w[166][6] = 5'b01111; w[166][7] = 5'b01111; w[166][8] = 5'b01111; w[166][9] = 5'b01111; w[166][10] = 5'b01111; w[166][11] = 5'b01111; w[166][12] = 5'b01111; w[166][13] = 5'b01111; w[166][14] = 5'b01111; w[166][15] = 5'b01111; w[166][16] = 5'b01111; w[166][17] = 5'b01111; w[166][18] = 5'b01111; w[166][19] = 5'b01111; w[166][20] = 5'b01111; w[166][21] = 5'b01111; w[166][22] = 5'b01111; w[166][23] = 5'b01111; w[166][24] = 5'b01111; w[166][25] = 5'b01111; w[166][26] = 5'b01111; w[166][27] = 5'b01111; w[166][28] = 5'b01111; w[166][29] = 5'b01111; w[166][30] = 5'b01111; w[166][31] = 5'b00000; w[166][32] = 5'b10000; w[166][33] = 5'b10000; w[166][34] = 5'b10000; w[166][35] = 5'b10000; w[166][36] = 5'b10000; w[166][37] = 5'b10000; w[166][38] = 5'b00000; w[166][39] = 5'b01111; w[166][40] = 5'b01111; w[166][41] = 5'b01111; w[166][42] = 5'b01111; w[166][43] = 5'b01111; w[166][44] = 5'b01111; w[166][45] = 5'b10000; w[166][46] = 5'b10000; w[166][47] = 5'b10000; w[166][48] = 5'b10000; w[166][49] = 5'b10000; w[166][50] = 5'b10000; w[166][51] = 5'b10000; w[166][52] = 5'b10000; w[166][53] = 5'b01111; w[166][54] = 5'b01111; w[166][55] = 5'b01111; w[166][56] = 5'b01111; w[166][57] = 5'b01111; w[166][58] = 5'b01111; w[166][59] = 5'b00000; w[166][60] = 5'b00000; w[166][61] = 5'b01111; w[166][62] = 5'b10000; w[166][63] = 5'b00000; w[166][64] = 5'b01111; w[166][65] = 5'b00000; w[166][66] = 5'b00000; w[166][67] = 5'b01111; w[166][68] = 5'b01111; w[166][69] = 5'b01111; w[166][70] = 5'b01111; w[166][71] = 5'b01111; w[166][72] = 5'b01111; w[166][73] = 5'b00000; w[166][74] = 5'b01111; w[166][75] = 5'b01111; w[166][76] = 5'b10000; w[166][77] = 5'b00000; w[166][78] = 5'b01111; w[166][79] = 5'b01111; w[166][80] = 5'b00000; w[166][81] = 5'b01111; w[166][82] = 5'b01111; w[166][83] = 5'b01111; w[166][84] = 5'b01111; w[166][85] = 5'b01111; w[166][86] = 5'b01111; w[166][87] = 5'b00000; w[166][88] = 5'b01111; w[166][89] = 5'b01111; w[166][90] = 5'b10000; w[166][91] = 5'b10000; w[166][92] = 5'b01111; w[166][93] = 5'b01111; w[166][94] = 5'b01111; w[166][95] = 5'b01111; w[166][96] = 5'b01111; w[166][97] = 5'b01111; w[166][98] = 5'b01111; w[166][99] = 5'b01111; w[166][100] = 5'b01111; w[166][101] = 5'b00000; w[166][102] = 5'b01111; w[166][103] = 5'b01111; w[166][104] = 5'b10000; w[166][105] = 5'b10000; w[166][106] = 5'b01111; w[166][107] = 5'b00000; w[166][108] = 5'b00000; w[166][109] = 5'b01111; w[166][110] = 5'b01111; w[166][111] = 5'b01111; w[166][112] = 5'b01111; w[166][113] = 5'b01111; w[166][114] = 5'b01111; w[166][115] = 5'b00000; w[166][116] = 5'b01111; w[166][117] = 5'b01111; w[166][118] = 5'b10000; w[166][119] = 5'b10000; w[166][120] = 5'b00000; w[166][121] = 5'b00000; w[166][122] = 5'b00000; w[166][123] = 5'b01111; w[166][124] = 5'b01111; w[166][125] = 5'b01111; w[166][126] = 5'b01111; w[166][127] = 5'b01111; w[166][128] = 5'b01111; w[166][129] = 5'b00000; w[166][130] = 5'b01111; w[166][131] = 5'b01111; w[166][132] = 5'b00000; w[166][133] = 5'b10000; w[166][134] = 5'b01111; w[166][135] = 5'b01111; w[166][136] = 5'b00000; w[166][137] = 5'b01111; w[166][138] = 5'b01111; w[166][139] = 5'b01111; w[166][140] = 5'b01111; w[166][141] = 5'b01111; w[166][142] = 5'b01111; w[166][143] = 5'b00000; w[166][144] = 5'b00000; w[166][145] = 5'b01111; w[166][146] = 5'b00000; w[166][147] = 5'b10000; w[166][148] = 5'b01111; w[166][149] = 5'b00000; w[166][150] = 5'b00000; w[166][151] = 5'b01111; w[166][152] = 5'b01111; w[166][153] = 5'b01111; w[166][154] = 5'b01111; w[166][155] = 5'b01111; w[166][156] = 5'b01111; w[166][157] = 5'b00000; w[166][158] = 5'b00000; w[166][159] = 5'b00000; w[166][160] = 5'b10000; w[166][161] = 5'b10000; w[166][162] = 5'b10000; w[166][163] = 5'b00000; w[166][164] = 5'b00000; w[166][165] = 5'b01111; w[166][166] = 5'b00000; w[166][167] = 5'b01111; w[166][168] = 5'b01111; w[166][169] = 5'b01111; w[166][170] = 5'b01111; w[166][171] = 5'b01111; w[166][172] = 5'b00000; w[166][173] = 5'b00000; w[166][174] = 5'b10000; w[166][175] = 5'b10000; w[166][176] = 5'b10000; w[166][177] = 5'b00000; w[166][178] = 5'b01111; w[166][179] = 5'b01111; w[166][180] = 5'b01111; w[166][181] = 5'b01111; w[166][182] = 5'b01111; w[166][183] = 5'b01111; w[166][184] = 5'b01111; w[166][185] = 5'b01111; w[166][186] = 5'b01111; w[166][187] = 5'b01111; w[166][188] = 5'b01111; w[166][189] = 5'b01111; w[166][190] = 5'b01111; w[166][191] = 5'b01111; w[166][192] = 5'b01111; w[166][193] = 5'b01111; w[166][194] = 5'b01111; w[166][195] = 5'b01111; w[166][196] = 5'b01111; w[166][197] = 5'b01111; w[166][198] = 5'b01111; w[166][199] = 5'b01111; w[166][200] = 5'b01111; w[166][201] = 5'b01111; w[166][202] = 5'b01111; w[166][203] = 5'b01111; w[166][204] = 5'b01111; w[166][205] = 5'b01111; w[166][206] = 5'b01111; w[166][207] = 5'b01111; w[166][208] = 5'b01111; w[166][209] = 5'b01111; 
w[167][0] = 5'b01111; w[167][1] = 5'b01111; w[167][2] = 5'b01111; w[167][3] = 5'b01111; w[167][4] = 5'b01111; w[167][5] = 5'b01111; w[167][6] = 5'b01111; w[167][7] = 5'b01111; w[167][8] = 5'b01111; w[167][9] = 5'b01111; w[167][10] = 5'b01111; w[167][11] = 5'b01111; w[167][12] = 5'b01111; w[167][13] = 5'b01111; w[167][14] = 5'b01111; w[167][15] = 5'b01111; w[167][16] = 5'b01111; w[167][17] = 5'b01111; w[167][18] = 5'b01111; w[167][19] = 5'b01111; w[167][20] = 5'b01111; w[167][21] = 5'b01111; w[167][22] = 5'b01111; w[167][23] = 5'b01111; w[167][24] = 5'b01111; w[167][25] = 5'b01111; w[167][26] = 5'b01111; w[167][27] = 5'b01111; w[167][28] = 5'b01111; w[167][29] = 5'b01111; w[167][30] = 5'b01111; w[167][31] = 5'b00000; w[167][32] = 5'b10000; w[167][33] = 5'b10000; w[167][34] = 5'b10000; w[167][35] = 5'b10000; w[167][36] = 5'b10000; w[167][37] = 5'b10000; w[167][38] = 5'b00000; w[167][39] = 5'b01111; w[167][40] = 5'b01111; w[167][41] = 5'b01111; w[167][42] = 5'b01111; w[167][43] = 5'b01111; w[167][44] = 5'b01111; w[167][45] = 5'b10000; w[167][46] = 5'b10000; w[167][47] = 5'b10000; w[167][48] = 5'b10000; w[167][49] = 5'b10000; w[167][50] = 5'b10000; w[167][51] = 5'b10000; w[167][52] = 5'b10000; w[167][53] = 5'b01111; w[167][54] = 5'b01111; w[167][55] = 5'b01111; w[167][56] = 5'b01111; w[167][57] = 5'b01111; w[167][58] = 5'b01111; w[167][59] = 5'b00000; w[167][60] = 5'b00000; w[167][61] = 5'b01111; w[167][62] = 5'b10000; w[167][63] = 5'b00000; w[167][64] = 5'b01111; w[167][65] = 5'b00000; w[167][66] = 5'b00000; w[167][67] = 5'b01111; w[167][68] = 5'b01111; w[167][69] = 5'b01111; w[167][70] = 5'b01111; w[167][71] = 5'b01111; w[167][72] = 5'b01111; w[167][73] = 5'b00000; w[167][74] = 5'b01111; w[167][75] = 5'b01111; w[167][76] = 5'b10000; w[167][77] = 5'b00000; w[167][78] = 5'b01111; w[167][79] = 5'b01111; w[167][80] = 5'b00000; w[167][81] = 5'b01111; w[167][82] = 5'b01111; w[167][83] = 5'b01111; w[167][84] = 5'b01111; w[167][85] = 5'b01111; w[167][86] = 5'b01111; w[167][87] = 5'b00000; w[167][88] = 5'b01111; w[167][89] = 5'b01111; w[167][90] = 5'b10000; w[167][91] = 5'b10000; w[167][92] = 5'b01111; w[167][93] = 5'b01111; w[167][94] = 5'b01111; w[167][95] = 5'b01111; w[167][96] = 5'b01111; w[167][97] = 5'b01111; w[167][98] = 5'b01111; w[167][99] = 5'b01111; w[167][100] = 5'b01111; w[167][101] = 5'b00000; w[167][102] = 5'b01111; w[167][103] = 5'b01111; w[167][104] = 5'b10000; w[167][105] = 5'b10000; w[167][106] = 5'b01111; w[167][107] = 5'b00000; w[167][108] = 5'b00000; w[167][109] = 5'b01111; w[167][110] = 5'b01111; w[167][111] = 5'b01111; w[167][112] = 5'b01111; w[167][113] = 5'b01111; w[167][114] = 5'b01111; w[167][115] = 5'b00000; w[167][116] = 5'b01111; w[167][117] = 5'b01111; w[167][118] = 5'b10000; w[167][119] = 5'b10000; w[167][120] = 5'b00000; w[167][121] = 5'b00000; w[167][122] = 5'b00000; w[167][123] = 5'b01111; w[167][124] = 5'b01111; w[167][125] = 5'b01111; w[167][126] = 5'b01111; w[167][127] = 5'b01111; w[167][128] = 5'b01111; w[167][129] = 5'b00000; w[167][130] = 5'b01111; w[167][131] = 5'b01111; w[167][132] = 5'b00000; w[167][133] = 5'b10000; w[167][134] = 5'b01111; w[167][135] = 5'b01111; w[167][136] = 5'b00000; w[167][137] = 5'b01111; w[167][138] = 5'b01111; w[167][139] = 5'b01111; w[167][140] = 5'b01111; w[167][141] = 5'b01111; w[167][142] = 5'b01111; w[167][143] = 5'b00000; w[167][144] = 5'b00000; w[167][145] = 5'b01111; w[167][146] = 5'b00000; w[167][147] = 5'b10000; w[167][148] = 5'b01111; w[167][149] = 5'b00000; w[167][150] = 5'b00000; w[167][151] = 5'b01111; w[167][152] = 5'b01111; w[167][153] = 5'b01111; w[167][154] = 5'b01111; w[167][155] = 5'b01111; w[167][156] = 5'b01111; w[167][157] = 5'b00000; w[167][158] = 5'b00000; w[167][159] = 5'b00000; w[167][160] = 5'b10000; w[167][161] = 5'b10000; w[167][162] = 5'b10000; w[167][163] = 5'b00000; w[167][164] = 5'b00000; w[167][165] = 5'b01111; w[167][166] = 5'b01111; w[167][167] = 5'b00000; w[167][168] = 5'b01111; w[167][169] = 5'b01111; w[167][170] = 5'b01111; w[167][171] = 5'b01111; w[167][172] = 5'b00000; w[167][173] = 5'b00000; w[167][174] = 5'b10000; w[167][175] = 5'b10000; w[167][176] = 5'b10000; w[167][177] = 5'b00000; w[167][178] = 5'b01111; w[167][179] = 5'b01111; w[167][180] = 5'b01111; w[167][181] = 5'b01111; w[167][182] = 5'b01111; w[167][183] = 5'b01111; w[167][184] = 5'b01111; w[167][185] = 5'b01111; w[167][186] = 5'b01111; w[167][187] = 5'b01111; w[167][188] = 5'b01111; w[167][189] = 5'b01111; w[167][190] = 5'b01111; w[167][191] = 5'b01111; w[167][192] = 5'b01111; w[167][193] = 5'b01111; w[167][194] = 5'b01111; w[167][195] = 5'b01111; w[167][196] = 5'b01111; w[167][197] = 5'b01111; w[167][198] = 5'b01111; w[167][199] = 5'b01111; w[167][200] = 5'b01111; w[167][201] = 5'b01111; w[167][202] = 5'b01111; w[167][203] = 5'b01111; w[167][204] = 5'b01111; w[167][205] = 5'b01111; w[167][206] = 5'b01111; w[167][207] = 5'b01111; w[167][208] = 5'b01111; w[167][209] = 5'b01111; 
w[168][0] = 5'b01111; w[168][1] = 5'b01111; w[168][2] = 5'b01111; w[168][3] = 5'b01111; w[168][4] = 5'b01111; w[168][5] = 5'b01111; w[168][6] = 5'b01111; w[168][7] = 5'b01111; w[168][8] = 5'b01111; w[168][9] = 5'b01111; w[168][10] = 5'b01111; w[168][11] = 5'b01111; w[168][12] = 5'b01111; w[168][13] = 5'b01111; w[168][14] = 5'b01111; w[168][15] = 5'b01111; w[168][16] = 5'b01111; w[168][17] = 5'b01111; w[168][18] = 5'b01111; w[168][19] = 5'b01111; w[168][20] = 5'b01111; w[168][21] = 5'b01111; w[168][22] = 5'b01111; w[168][23] = 5'b01111; w[168][24] = 5'b01111; w[168][25] = 5'b01111; w[168][26] = 5'b01111; w[168][27] = 5'b01111; w[168][28] = 5'b01111; w[168][29] = 5'b01111; w[168][30] = 5'b01111; w[168][31] = 5'b00000; w[168][32] = 5'b10000; w[168][33] = 5'b10000; w[168][34] = 5'b10000; w[168][35] = 5'b10000; w[168][36] = 5'b10000; w[168][37] = 5'b10000; w[168][38] = 5'b00000; w[168][39] = 5'b01111; w[168][40] = 5'b01111; w[168][41] = 5'b01111; w[168][42] = 5'b01111; w[168][43] = 5'b01111; w[168][44] = 5'b01111; w[168][45] = 5'b10000; w[168][46] = 5'b10000; w[168][47] = 5'b10000; w[168][48] = 5'b10000; w[168][49] = 5'b10000; w[168][50] = 5'b10000; w[168][51] = 5'b10000; w[168][52] = 5'b10000; w[168][53] = 5'b01111; w[168][54] = 5'b01111; w[168][55] = 5'b01111; w[168][56] = 5'b01111; w[168][57] = 5'b01111; w[168][58] = 5'b01111; w[168][59] = 5'b00000; w[168][60] = 5'b00000; w[168][61] = 5'b01111; w[168][62] = 5'b10000; w[168][63] = 5'b00000; w[168][64] = 5'b01111; w[168][65] = 5'b00000; w[168][66] = 5'b00000; w[168][67] = 5'b01111; w[168][68] = 5'b01111; w[168][69] = 5'b01111; w[168][70] = 5'b01111; w[168][71] = 5'b01111; w[168][72] = 5'b01111; w[168][73] = 5'b00000; w[168][74] = 5'b01111; w[168][75] = 5'b01111; w[168][76] = 5'b10000; w[168][77] = 5'b00000; w[168][78] = 5'b01111; w[168][79] = 5'b01111; w[168][80] = 5'b00000; w[168][81] = 5'b01111; w[168][82] = 5'b01111; w[168][83] = 5'b01111; w[168][84] = 5'b01111; w[168][85] = 5'b01111; w[168][86] = 5'b01111; w[168][87] = 5'b00000; w[168][88] = 5'b01111; w[168][89] = 5'b01111; w[168][90] = 5'b10000; w[168][91] = 5'b10000; w[168][92] = 5'b01111; w[168][93] = 5'b01111; w[168][94] = 5'b01111; w[168][95] = 5'b01111; w[168][96] = 5'b01111; w[168][97] = 5'b01111; w[168][98] = 5'b01111; w[168][99] = 5'b01111; w[168][100] = 5'b01111; w[168][101] = 5'b00000; w[168][102] = 5'b01111; w[168][103] = 5'b01111; w[168][104] = 5'b10000; w[168][105] = 5'b10000; w[168][106] = 5'b01111; w[168][107] = 5'b00000; w[168][108] = 5'b00000; w[168][109] = 5'b01111; w[168][110] = 5'b01111; w[168][111] = 5'b01111; w[168][112] = 5'b01111; w[168][113] = 5'b01111; w[168][114] = 5'b01111; w[168][115] = 5'b00000; w[168][116] = 5'b01111; w[168][117] = 5'b01111; w[168][118] = 5'b10000; w[168][119] = 5'b10000; w[168][120] = 5'b00000; w[168][121] = 5'b00000; w[168][122] = 5'b00000; w[168][123] = 5'b01111; w[168][124] = 5'b01111; w[168][125] = 5'b01111; w[168][126] = 5'b01111; w[168][127] = 5'b01111; w[168][128] = 5'b01111; w[168][129] = 5'b00000; w[168][130] = 5'b01111; w[168][131] = 5'b01111; w[168][132] = 5'b00000; w[168][133] = 5'b10000; w[168][134] = 5'b01111; w[168][135] = 5'b01111; w[168][136] = 5'b00000; w[168][137] = 5'b01111; w[168][138] = 5'b01111; w[168][139] = 5'b01111; w[168][140] = 5'b01111; w[168][141] = 5'b01111; w[168][142] = 5'b01111; w[168][143] = 5'b00000; w[168][144] = 5'b00000; w[168][145] = 5'b01111; w[168][146] = 5'b00000; w[168][147] = 5'b10000; w[168][148] = 5'b01111; w[168][149] = 5'b00000; w[168][150] = 5'b00000; w[168][151] = 5'b01111; w[168][152] = 5'b01111; w[168][153] = 5'b01111; w[168][154] = 5'b01111; w[168][155] = 5'b01111; w[168][156] = 5'b01111; w[168][157] = 5'b00000; w[168][158] = 5'b00000; w[168][159] = 5'b00000; w[168][160] = 5'b10000; w[168][161] = 5'b10000; w[168][162] = 5'b10000; w[168][163] = 5'b00000; w[168][164] = 5'b00000; w[168][165] = 5'b01111; w[168][166] = 5'b01111; w[168][167] = 5'b01111; w[168][168] = 5'b00000; w[168][169] = 5'b01111; w[168][170] = 5'b01111; w[168][171] = 5'b01111; w[168][172] = 5'b00000; w[168][173] = 5'b00000; w[168][174] = 5'b10000; w[168][175] = 5'b10000; w[168][176] = 5'b10000; w[168][177] = 5'b00000; w[168][178] = 5'b01111; w[168][179] = 5'b01111; w[168][180] = 5'b01111; w[168][181] = 5'b01111; w[168][182] = 5'b01111; w[168][183] = 5'b01111; w[168][184] = 5'b01111; w[168][185] = 5'b01111; w[168][186] = 5'b01111; w[168][187] = 5'b01111; w[168][188] = 5'b01111; w[168][189] = 5'b01111; w[168][190] = 5'b01111; w[168][191] = 5'b01111; w[168][192] = 5'b01111; w[168][193] = 5'b01111; w[168][194] = 5'b01111; w[168][195] = 5'b01111; w[168][196] = 5'b01111; w[168][197] = 5'b01111; w[168][198] = 5'b01111; w[168][199] = 5'b01111; w[168][200] = 5'b01111; w[168][201] = 5'b01111; w[168][202] = 5'b01111; w[168][203] = 5'b01111; w[168][204] = 5'b01111; w[168][205] = 5'b01111; w[168][206] = 5'b01111; w[168][207] = 5'b01111; w[168][208] = 5'b01111; w[168][209] = 5'b01111; 
w[169][0] = 5'b01111; w[169][1] = 5'b01111; w[169][2] = 5'b01111; w[169][3] = 5'b01111; w[169][4] = 5'b01111; w[169][5] = 5'b01111; w[169][6] = 5'b01111; w[169][7] = 5'b01111; w[169][8] = 5'b01111; w[169][9] = 5'b01111; w[169][10] = 5'b01111; w[169][11] = 5'b01111; w[169][12] = 5'b01111; w[169][13] = 5'b01111; w[169][14] = 5'b01111; w[169][15] = 5'b01111; w[169][16] = 5'b01111; w[169][17] = 5'b01111; w[169][18] = 5'b01111; w[169][19] = 5'b01111; w[169][20] = 5'b01111; w[169][21] = 5'b01111; w[169][22] = 5'b01111; w[169][23] = 5'b01111; w[169][24] = 5'b01111; w[169][25] = 5'b01111; w[169][26] = 5'b01111; w[169][27] = 5'b01111; w[169][28] = 5'b01111; w[169][29] = 5'b01111; w[169][30] = 5'b01111; w[169][31] = 5'b00000; w[169][32] = 5'b10000; w[169][33] = 5'b10000; w[169][34] = 5'b10000; w[169][35] = 5'b10000; w[169][36] = 5'b10000; w[169][37] = 5'b10000; w[169][38] = 5'b00000; w[169][39] = 5'b01111; w[169][40] = 5'b01111; w[169][41] = 5'b01111; w[169][42] = 5'b01111; w[169][43] = 5'b01111; w[169][44] = 5'b01111; w[169][45] = 5'b10000; w[169][46] = 5'b10000; w[169][47] = 5'b10000; w[169][48] = 5'b10000; w[169][49] = 5'b10000; w[169][50] = 5'b10000; w[169][51] = 5'b10000; w[169][52] = 5'b10000; w[169][53] = 5'b01111; w[169][54] = 5'b01111; w[169][55] = 5'b01111; w[169][56] = 5'b01111; w[169][57] = 5'b01111; w[169][58] = 5'b01111; w[169][59] = 5'b00000; w[169][60] = 5'b00000; w[169][61] = 5'b01111; w[169][62] = 5'b10000; w[169][63] = 5'b00000; w[169][64] = 5'b01111; w[169][65] = 5'b00000; w[169][66] = 5'b00000; w[169][67] = 5'b01111; w[169][68] = 5'b01111; w[169][69] = 5'b01111; w[169][70] = 5'b01111; w[169][71] = 5'b01111; w[169][72] = 5'b01111; w[169][73] = 5'b00000; w[169][74] = 5'b01111; w[169][75] = 5'b01111; w[169][76] = 5'b10000; w[169][77] = 5'b00000; w[169][78] = 5'b01111; w[169][79] = 5'b01111; w[169][80] = 5'b00000; w[169][81] = 5'b01111; w[169][82] = 5'b01111; w[169][83] = 5'b01111; w[169][84] = 5'b01111; w[169][85] = 5'b01111; w[169][86] = 5'b01111; w[169][87] = 5'b00000; w[169][88] = 5'b01111; w[169][89] = 5'b01111; w[169][90] = 5'b10000; w[169][91] = 5'b10000; w[169][92] = 5'b01111; w[169][93] = 5'b01111; w[169][94] = 5'b01111; w[169][95] = 5'b01111; w[169][96] = 5'b01111; w[169][97] = 5'b01111; w[169][98] = 5'b01111; w[169][99] = 5'b01111; w[169][100] = 5'b01111; w[169][101] = 5'b00000; w[169][102] = 5'b01111; w[169][103] = 5'b01111; w[169][104] = 5'b10000; w[169][105] = 5'b10000; w[169][106] = 5'b01111; w[169][107] = 5'b00000; w[169][108] = 5'b00000; w[169][109] = 5'b01111; w[169][110] = 5'b01111; w[169][111] = 5'b01111; w[169][112] = 5'b01111; w[169][113] = 5'b01111; w[169][114] = 5'b01111; w[169][115] = 5'b00000; w[169][116] = 5'b01111; w[169][117] = 5'b01111; w[169][118] = 5'b10000; w[169][119] = 5'b10000; w[169][120] = 5'b00000; w[169][121] = 5'b00000; w[169][122] = 5'b00000; w[169][123] = 5'b01111; w[169][124] = 5'b01111; w[169][125] = 5'b01111; w[169][126] = 5'b01111; w[169][127] = 5'b01111; w[169][128] = 5'b01111; w[169][129] = 5'b00000; w[169][130] = 5'b01111; w[169][131] = 5'b01111; w[169][132] = 5'b00000; w[169][133] = 5'b10000; w[169][134] = 5'b01111; w[169][135] = 5'b01111; w[169][136] = 5'b00000; w[169][137] = 5'b01111; w[169][138] = 5'b01111; w[169][139] = 5'b01111; w[169][140] = 5'b01111; w[169][141] = 5'b01111; w[169][142] = 5'b01111; w[169][143] = 5'b00000; w[169][144] = 5'b00000; w[169][145] = 5'b01111; w[169][146] = 5'b00000; w[169][147] = 5'b10000; w[169][148] = 5'b01111; w[169][149] = 5'b00000; w[169][150] = 5'b00000; w[169][151] = 5'b01111; w[169][152] = 5'b01111; w[169][153] = 5'b01111; w[169][154] = 5'b01111; w[169][155] = 5'b01111; w[169][156] = 5'b01111; w[169][157] = 5'b00000; w[169][158] = 5'b00000; w[169][159] = 5'b00000; w[169][160] = 5'b10000; w[169][161] = 5'b10000; w[169][162] = 5'b10000; w[169][163] = 5'b00000; w[169][164] = 5'b00000; w[169][165] = 5'b01111; w[169][166] = 5'b01111; w[169][167] = 5'b01111; w[169][168] = 5'b01111; w[169][169] = 5'b00000; w[169][170] = 5'b01111; w[169][171] = 5'b01111; w[169][172] = 5'b00000; w[169][173] = 5'b00000; w[169][174] = 5'b10000; w[169][175] = 5'b10000; w[169][176] = 5'b10000; w[169][177] = 5'b00000; w[169][178] = 5'b01111; w[169][179] = 5'b01111; w[169][180] = 5'b01111; w[169][181] = 5'b01111; w[169][182] = 5'b01111; w[169][183] = 5'b01111; w[169][184] = 5'b01111; w[169][185] = 5'b01111; w[169][186] = 5'b01111; w[169][187] = 5'b01111; w[169][188] = 5'b01111; w[169][189] = 5'b01111; w[169][190] = 5'b01111; w[169][191] = 5'b01111; w[169][192] = 5'b01111; w[169][193] = 5'b01111; w[169][194] = 5'b01111; w[169][195] = 5'b01111; w[169][196] = 5'b01111; w[169][197] = 5'b01111; w[169][198] = 5'b01111; w[169][199] = 5'b01111; w[169][200] = 5'b01111; w[169][201] = 5'b01111; w[169][202] = 5'b01111; w[169][203] = 5'b01111; w[169][204] = 5'b01111; w[169][205] = 5'b01111; w[169][206] = 5'b01111; w[169][207] = 5'b01111; w[169][208] = 5'b01111; w[169][209] = 5'b01111; 
w[170][0] = 5'b01111; w[170][1] = 5'b01111; w[170][2] = 5'b01111; w[170][3] = 5'b01111; w[170][4] = 5'b01111; w[170][5] = 5'b01111; w[170][6] = 5'b01111; w[170][7] = 5'b01111; w[170][8] = 5'b01111; w[170][9] = 5'b01111; w[170][10] = 5'b01111; w[170][11] = 5'b01111; w[170][12] = 5'b01111; w[170][13] = 5'b01111; w[170][14] = 5'b01111; w[170][15] = 5'b01111; w[170][16] = 5'b01111; w[170][17] = 5'b01111; w[170][18] = 5'b01111; w[170][19] = 5'b01111; w[170][20] = 5'b01111; w[170][21] = 5'b01111; w[170][22] = 5'b01111; w[170][23] = 5'b01111; w[170][24] = 5'b01111; w[170][25] = 5'b01111; w[170][26] = 5'b01111; w[170][27] = 5'b01111; w[170][28] = 5'b01111; w[170][29] = 5'b01111; w[170][30] = 5'b01111; w[170][31] = 5'b00000; w[170][32] = 5'b10000; w[170][33] = 5'b10000; w[170][34] = 5'b10000; w[170][35] = 5'b10000; w[170][36] = 5'b10000; w[170][37] = 5'b10000; w[170][38] = 5'b00000; w[170][39] = 5'b01111; w[170][40] = 5'b01111; w[170][41] = 5'b01111; w[170][42] = 5'b01111; w[170][43] = 5'b01111; w[170][44] = 5'b01111; w[170][45] = 5'b10000; w[170][46] = 5'b10000; w[170][47] = 5'b10000; w[170][48] = 5'b10000; w[170][49] = 5'b10000; w[170][50] = 5'b10000; w[170][51] = 5'b10000; w[170][52] = 5'b10000; w[170][53] = 5'b01111; w[170][54] = 5'b01111; w[170][55] = 5'b01111; w[170][56] = 5'b01111; w[170][57] = 5'b01111; w[170][58] = 5'b01111; w[170][59] = 5'b00000; w[170][60] = 5'b00000; w[170][61] = 5'b01111; w[170][62] = 5'b10000; w[170][63] = 5'b00000; w[170][64] = 5'b01111; w[170][65] = 5'b00000; w[170][66] = 5'b00000; w[170][67] = 5'b01111; w[170][68] = 5'b01111; w[170][69] = 5'b01111; w[170][70] = 5'b01111; w[170][71] = 5'b01111; w[170][72] = 5'b01111; w[170][73] = 5'b00000; w[170][74] = 5'b01111; w[170][75] = 5'b01111; w[170][76] = 5'b10000; w[170][77] = 5'b00000; w[170][78] = 5'b01111; w[170][79] = 5'b01111; w[170][80] = 5'b00000; w[170][81] = 5'b01111; w[170][82] = 5'b01111; w[170][83] = 5'b01111; w[170][84] = 5'b01111; w[170][85] = 5'b01111; w[170][86] = 5'b01111; w[170][87] = 5'b00000; w[170][88] = 5'b01111; w[170][89] = 5'b01111; w[170][90] = 5'b10000; w[170][91] = 5'b10000; w[170][92] = 5'b01111; w[170][93] = 5'b01111; w[170][94] = 5'b01111; w[170][95] = 5'b01111; w[170][96] = 5'b01111; w[170][97] = 5'b01111; w[170][98] = 5'b01111; w[170][99] = 5'b01111; w[170][100] = 5'b01111; w[170][101] = 5'b00000; w[170][102] = 5'b01111; w[170][103] = 5'b01111; w[170][104] = 5'b10000; w[170][105] = 5'b10000; w[170][106] = 5'b01111; w[170][107] = 5'b00000; w[170][108] = 5'b00000; w[170][109] = 5'b01111; w[170][110] = 5'b01111; w[170][111] = 5'b01111; w[170][112] = 5'b01111; w[170][113] = 5'b01111; w[170][114] = 5'b01111; w[170][115] = 5'b00000; w[170][116] = 5'b01111; w[170][117] = 5'b01111; w[170][118] = 5'b10000; w[170][119] = 5'b10000; w[170][120] = 5'b00000; w[170][121] = 5'b00000; w[170][122] = 5'b00000; w[170][123] = 5'b01111; w[170][124] = 5'b01111; w[170][125] = 5'b01111; w[170][126] = 5'b01111; w[170][127] = 5'b01111; w[170][128] = 5'b01111; w[170][129] = 5'b00000; w[170][130] = 5'b01111; w[170][131] = 5'b01111; w[170][132] = 5'b00000; w[170][133] = 5'b10000; w[170][134] = 5'b01111; w[170][135] = 5'b01111; w[170][136] = 5'b00000; w[170][137] = 5'b01111; w[170][138] = 5'b01111; w[170][139] = 5'b01111; w[170][140] = 5'b01111; w[170][141] = 5'b01111; w[170][142] = 5'b01111; w[170][143] = 5'b00000; w[170][144] = 5'b00000; w[170][145] = 5'b01111; w[170][146] = 5'b00000; w[170][147] = 5'b10000; w[170][148] = 5'b01111; w[170][149] = 5'b00000; w[170][150] = 5'b00000; w[170][151] = 5'b01111; w[170][152] = 5'b01111; w[170][153] = 5'b01111; w[170][154] = 5'b01111; w[170][155] = 5'b01111; w[170][156] = 5'b01111; w[170][157] = 5'b00000; w[170][158] = 5'b00000; w[170][159] = 5'b00000; w[170][160] = 5'b10000; w[170][161] = 5'b10000; w[170][162] = 5'b10000; w[170][163] = 5'b00000; w[170][164] = 5'b00000; w[170][165] = 5'b01111; w[170][166] = 5'b01111; w[170][167] = 5'b01111; w[170][168] = 5'b01111; w[170][169] = 5'b01111; w[170][170] = 5'b00000; w[170][171] = 5'b01111; w[170][172] = 5'b00000; w[170][173] = 5'b00000; w[170][174] = 5'b10000; w[170][175] = 5'b10000; w[170][176] = 5'b10000; w[170][177] = 5'b00000; w[170][178] = 5'b01111; w[170][179] = 5'b01111; w[170][180] = 5'b01111; w[170][181] = 5'b01111; w[170][182] = 5'b01111; w[170][183] = 5'b01111; w[170][184] = 5'b01111; w[170][185] = 5'b01111; w[170][186] = 5'b01111; w[170][187] = 5'b01111; w[170][188] = 5'b01111; w[170][189] = 5'b01111; w[170][190] = 5'b01111; w[170][191] = 5'b01111; w[170][192] = 5'b01111; w[170][193] = 5'b01111; w[170][194] = 5'b01111; w[170][195] = 5'b01111; w[170][196] = 5'b01111; w[170][197] = 5'b01111; w[170][198] = 5'b01111; w[170][199] = 5'b01111; w[170][200] = 5'b01111; w[170][201] = 5'b01111; w[170][202] = 5'b01111; w[170][203] = 5'b01111; w[170][204] = 5'b01111; w[170][205] = 5'b01111; w[170][206] = 5'b01111; w[170][207] = 5'b01111; w[170][208] = 5'b01111; w[170][209] = 5'b01111; 
w[171][0] = 5'b01111; w[171][1] = 5'b01111; w[171][2] = 5'b01111; w[171][3] = 5'b01111; w[171][4] = 5'b01111; w[171][5] = 5'b01111; w[171][6] = 5'b01111; w[171][7] = 5'b01111; w[171][8] = 5'b01111; w[171][9] = 5'b01111; w[171][10] = 5'b01111; w[171][11] = 5'b01111; w[171][12] = 5'b01111; w[171][13] = 5'b01111; w[171][14] = 5'b01111; w[171][15] = 5'b01111; w[171][16] = 5'b01111; w[171][17] = 5'b01111; w[171][18] = 5'b01111; w[171][19] = 5'b01111; w[171][20] = 5'b01111; w[171][21] = 5'b01111; w[171][22] = 5'b01111; w[171][23] = 5'b01111; w[171][24] = 5'b01111; w[171][25] = 5'b01111; w[171][26] = 5'b01111; w[171][27] = 5'b01111; w[171][28] = 5'b01111; w[171][29] = 5'b01111; w[171][30] = 5'b00000; w[171][31] = 5'b01111; w[171][32] = 5'b00000; w[171][33] = 5'b10000; w[171][34] = 5'b10000; w[171][35] = 5'b10000; w[171][36] = 5'b10000; w[171][37] = 5'b00000; w[171][38] = 5'b01111; w[171][39] = 5'b00000; w[171][40] = 5'b01111; w[171][41] = 5'b01111; w[171][42] = 5'b01111; w[171][43] = 5'b01111; w[171][44] = 5'b00000; w[171][45] = 5'b00000; w[171][46] = 5'b00000; w[171][47] = 5'b10000; w[171][48] = 5'b10000; w[171][49] = 5'b10000; w[171][50] = 5'b10000; w[171][51] = 5'b00000; w[171][52] = 5'b00000; w[171][53] = 5'b00000; w[171][54] = 5'b01111; w[171][55] = 5'b01111; w[171][56] = 5'b01111; w[171][57] = 5'b01111; w[171][58] = 5'b00000; w[171][59] = 5'b01111; w[171][60] = 5'b01111; w[171][61] = 5'b01111; w[171][62] = 5'b00000; w[171][63] = 5'b10000; w[171][64] = 5'b01111; w[171][65] = 5'b01111; w[171][66] = 5'b01111; w[171][67] = 5'b00000; w[171][68] = 5'b01111; w[171][69] = 5'b01111; w[171][70] = 5'b01111; w[171][71] = 5'b01111; w[171][72] = 5'b00000; w[171][73] = 5'b01111; w[171][74] = 5'b01111; w[171][75] = 5'b01111; w[171][76] = 5'b00000; w[171][77] = 5'b10000; w[171][78] = 5'b01111; w[171][79] = 5'b01111; w[171][80] = 5'b01111; w[171][81] = 5'b00000; w[171][82] = 5'b01111; w[171][83] = 5'b01111; w[171][84] = 5'b01111; w[171][85] = 5'b01111; w[171][86] = 5'b00000; w[171][87] = 5'b01111; w[171][88] = 5'b01111; w[171][89] = 5'b01111; w[171][90] = 5'b00000; w[171][91] = 5'b00000; w[171][92] = 5'b01111; w[171][93] = 5'b01111; w[171][94] = 5'b01111; w[171][95] = 5'b01111; w[171][96] = 5'b01111; w[171][97] = 5'b01111; w[171][98] = 5'b01111; w[171][99] = 5'b01111; w[171][100] = 5'b00000; w[171][101] = 5'b01111; w[171][102] = 5'b01111; w[171][103] = 5'b01111; w[171][104] = 5'b00000; w[171][105] = 5'b00000; w[171][106] = 5'b00000; w[171][107] = 5'b01111; w[171][108] = 5'b01111; w[171][109] = 5'b00000; w[171][110] = 5'b01111; w[171][111] = 5'b01111; w[171][112] = 5'b01111; w[171][113] = 5'b01111; w[171][114] = 5'b00000; w[171][115] = 5'b01111; w[171][116] = 5'b01111; w[171][117] = 5'b01111; w[171][118] = 5'b00000; w[171][119] = 5'b00000; w[171][120] = 5'b01111; w[171][121] = 5'b01111; w[171][122] = 5'b01111; w[171][123] = 5'b00000; w[171][124] = 5'b01111; w[171][125] = 5'b01111; w[171][126] = 5'b01111; w[171][127] = 5'b01111; w[171][128] = 5'b00000; w[171][129] = 5'b01111; w[171][130] = 5'b01111; w[171][131] = 5'b01111; w[171][132] = 5'b10000; w[171][133] = 5'b00000; w[171][134] = 5'b01111; w[171][135] = 5'b01111; w[171][136] = 5'b01111; w[171][137] = 5'b00000; w[171][138] = 5'b01111; w[171][139] = 5'b01111; w[171][140] = 5'b01111; w[171][141] = 5'b01111; w[171][142] = 5'b00000; w[171][143] = 5'b01111; w[171][144] = 5'b01111; w[171][145] = 5'b01111; w[171][146] = 5'b10000; w[171][147] = 5'b00000; w[171][148] = 5'b01111; w[171][149] = 5'b01111; w[171][150] = 5'b01111; w[171][151] = 5'b00000; w[171][152] = 5'b01111; w[171][153] = 5'b01111; w[171][154] = 5'b01111; w[171][155] = 5'b01111; w[171][156] = 5'b01111; w[171][157] = 5'b01111; w[171][158] = 5'b01111; w[171][159] = 5'b10000; w[171][160] = 5'b10000; w[171][161] = 5'b10000; w[171][162] = 5'b00000; w[171][163] = 5'b01111; w[171][164] = 5'b01111; w[171][165] = 5'b01111; w[171][166] = 5'b01111; w[171][167] = 5'b01111; w[171][168] = 5'b01111; w[171][169] = 5'b01111; w[171][170] = 5'b01111; w[171][171] = 5'b00000; w[171][172] = 5'b01111; w[171][173] = 5'b10000; w[171][174] = 5'b10000; w[171][175] = 5'b10000; w[171][176] = 5'b00000; w[171][177] = 5'b01111; w[171][178] = 5'b01111; w[171][179] = 5'b01111; w[171][180] = 5'b01111; w[171][181] = 5'b01111; w[171][182] = 5'b01111; w[171][183] = 5'b01111; w[171][184] = 5'b01111; w[171][185] = 5'b01111; w[171][186] = 5'b01111; w[171][187] = 5'b01111; w[171][188] = 5'b01111; w[171][189] = 5'b01111; w[171][190] = 5'b01111; w[171][191] = 5'b01111; w[171][192] = 5'b01111; w[171][193] = 5'b01111; w[171][194] = 5'b01111; w[171][195] = 5'b01111; w[171][196] = 5'b01111; w[171][197] = 5'b01111; w[171][198] = 5'b01111; w[171][199] = 5'b01111; w[171][200] = 5'b01111; w[171][201] = 5'b01111; w[171][202] = 5'b01111; w[171][203] = 5'b01111; w[171][204] = 5'b01111; w[171][205] = 5'b01111; w[171][206] = 5'b01111; w[171][207] = 5'b01111; w[171][208] = 5'b01111; w[171][209] = 5'b01111; 
w[172][0] = 5'b00000; w[172][1] = 5'b00000; w[172][2] = 5'b00000; w[172][3] = 5'b00000; w[172][4] = 5'b00000; w[172][5] = 5'b00000; w[172][6] = 5'b00000; w[172][7] = 5'b00000; w[172][8] = 5'b00000; w[172][9] = 5'b00000; w[172][10] = 5'b00000; w[172][11] = 5'b00000; w[172][12] = 5'b00000; w[172][13] = 5'b00000; w[172][14] = 5'b00000; w[172][15] = 5'b00000; w[172][16] = 5'b00000; w[172][17] = 5'b00000; w[172][18] = 5'b00000; w[172][19] = 5'b00000; w[172][20] = 5'b00000; w[172][21] = 5'b00000; w[172][22] = 5'b00000; w[172][23] = 5'b00000; w[172][24] = 5'b00000; w[172][25] = 5'b00000; w[172][26] = 5'b00000; w[172][27] = 5'b00000; w[172][28] = 5'b00000; w[172][29] = 5'b00000; w[172][30] = 5'b10000; w[172][31] = 5'b00000; w[172][32] = 5'b01111; w[172][33] = 5'b00000; w[172][34] = 5'b10000; w[172][35] = 5'b10000; w[172][36] = 5'b10000; w[172][37] = 5'b01111; w[172][38] = 5'b00000; w[172][39] = 5'b10000; w[172][40] = 5'b00000; w[172][41] = 5'b00000; w[172][42] = 5'b00000; w[172][43] = 5'b00000; w[172][44] = 5'b10000; w[172][45] = 5'b01111; w[172][46] = 5'b01111; w[172][47] = 5'b00000; w[172][48] = 5'b10000; w[172][49] = 5'b10000; w[172][50] = 5'b10000; w[172][51] = 5'b01111; w[172][52] = 5'b01111; w[172][53] = 5'b10000; w[172][54] = 5'b00000; w[172][55] = 5'b00000; w[172][56] = 5'b00000; w[172][57] = 5'b00000; w[172][58] = 5'b01111; w[172][59] = 5'b01111; w[172][60] = 5'b01111; w[172][61] = 5'b01111; w[172][62] = 5'b10000; w[172][63] = 5'b10000; w[172][64] = 5'b00000; w[172][65] = 5'b01111; w[172][66] = 5'b01111; w[172][67] = 5'b01111; w[172][68] = 5'b00000; w[172][69] = 5'b00000; w[172][70] = 5'b00000; w[172][71] = 5'b00000; w[172][72] = 5'b01111; w[172][73] = 5'b01111; w[172][74] = 5'b01111; w[172][75] = 5'b01111; w[172][76] = 5'b10000; w[172][77] = 5'b10000; w[172][78] = 5'b00000; w[172][79] = 5'b01111; w[172][80] = 5'b01111; w[172][81] = 5'b01111; w[172][82] = 5'b00000; w[172][83] = 5'b00000; w[172][84] = 5'b00000; w[172][85] = 5'b00000; w[172][86] = 5'b01111; w[172][87] = 5'b01111; w[172][88] = 5'b01111; w[172][89] = 5'b01111; w[172][90] = 5'b10000; w[172][91] = 5'b10000; w[172][92] = 5'b00000; w[172][93] = 5'b01111; w[172][94] = 5'b01111; w[172][95] = 5'b00000; w[172][96] = 5'b00000; w[172][97] = 5'b00000; w[172][98] = 5'b00000; w[172][99] = 5'b00000; w[172][100] = 5'b01111; w[172][101] = 5'b01111; w[172][102] = 5'b01111; w[172][103] = 5'b00000; w[172][104] = 5'b10000; w[172][105] = 5'b10000; w[172][106] = 5'b01111; w[172][107] = 5'b01111; w[172][108] = 5'b01111; w[172][109] = 5'b01111; w[172][110] = 5'b00000; w[172][111] = 5'b00000; w[172][112] = 5'b00000; w[172][113] = 5'b00000; w[172][114] = 5'b01111; w[172][115] = 5'b01111; w[172][116] = 5'b01111; w[172][117] = 5'b00000; w[172][118] = 5'b10000; w[172][119] = 5'b10000; w[172][120] = 5'b01111; w[172][121] = 5'b01111; w[172][122] = 5'b01111; w[172][123] = 5'b01111; w[172][124] = 5'b00000; w[172][125] = 5'b00000; w[172][126] = 5'b00000; w[172][127] = 5'b00000; w[172][128] = 5'b01111; w[172][129] = 5'b01111; w[172][130] = 5'b01111; w[172][131] = 5'b00000; w[172][132] = 5'b10000; w[172][133] = 5'b10000; w[172][134] = 5'b01111; w[172][135] = 5'b01111; w[172][136] = 5'b01111; w[172][137] = 5'b01111; w[172][138] = 5'b00000; w[172][139] = 5'b00000; w[172][140] = 5'b00000; w[172][141] = 5'b00000; w[172][142] = 5'b01111; w[172][143] = 5'b01111; w[172][144] = 5'b01111; w[172][145] = 5'b00000; w[172][146] = 5'b10000; w[172][147] = 5'b10000; w[172][148] = 5'b01111; w[172][149] = 5'b01111; w[172][150] = 5'b01111; w[172][151] = 5'b01111; w[172][152] = 5'b00000; w[172][153] = 5'b00000; w[172][154] = 5'b00000; w[172][155] = 5'b00000; w[172][156] = 5'b00000; w[172][157] = 5'b01111; w[172][158] = 5'b01111; w[172][159] = 5'b00000; w[172][160] = 5'b10000; w[172][161] = 5'b10000; w[172][162] = 5'b01111; w[172][163] = 5'b01111; w[172][164] = 5'b01111; w[172][165] = 5'b00000; w[172][166] = 5'b00000; w[172][167] = 5'b00000; w[172][168] = 5'b00000; w[172][169] = 5'b00000; w[172][170] = 5'b00000; w[172][171] = 5'b01111; w[172][172] = 5'b00000; w[172][173] = 5'b00000; w[172][174] = 5'b10000; w[172][175] = 5'b10000; w[172][176] = 5'b01111; w[172][177] = 5'b01111; w[172][178] = 5'b01111; w[172][179] = 5'b00000; w[172][180] = 5'b00000; w[172][181] = 5'b00000; w[172][182] = 5'b00000; w[172][183] = 5'b00000; w[172][184] = 5'b00000; w[172][185] = 5'b00000; w[172][186] = 5'b00000; w[172][187] = 5'b00000; w[172][188] = 5'b00000; w[172][189] = 5'b00000; w[172][190] = 5'b00000; w[172][191] = 5'b00000; w[172][192] = 5'b00000; w[172][193] = 5'b00000; w[172][194] = 5'b00000; w[172][195] = 5'b00000; w[172][196] = 5'b00000; w[172][197] = 5'b00000; w[172][198] = 5'b00000; w[172][199] = 5'b00000; w[172][200] = 5'b00000; w[172][201] = 5'b00000; w[172][202] = 5'b00000; w[172][203] = 5'b00000; w[172][204] = 5'b00000; w[172][205] = 5'b00000; w[172][206] = 5'b00000; w[172][207] = 5'b00000; w[172][208] = 5'b00000; w[172][209] = 5'b00000; 
w[173][0] = 5'b00000; w[173][1] = 5'b00000; w[173][2] = 5'b00000; w[173][3] = 5'b00000; w[173][4] = 5'b00000; w[173][5] = 5'b00000; w[173][6] = 5'b00000; w[173][7] = 5'b00000; w[173][8] = 5'b00000; w[173][9] = 5'b00000; w[173][10] = 5'b00000; w[173][11] = 5'b00000; w[173][12] = 5'b00000; w[173][13] = 5'b00000; w[173][14] = 5'b00000; w[173][15] = 5'b00000; w[173][16] = 5'b00000; w[173][17] = 5'b00000; w[173][18] = 5'b00000; w[173][19] = 5'b00000; w[173][20] = 5'b00000; w[173][21] = 5'b00000; w[173][22] = 5'b00000; w[173][23] = 5'b00000; w[173][24] = 5'b00000; w[173][25] = 5'b00000; w[173][26] = 5'b00000; w[173][27] = 5'b00000; w[173][28] = 5'b00000; w[173][29] = 5'b00000; w[173][30] = 5'b10000; w[173][31] = 5'b10000; w[173][32] = 5'b10000; w[173][33] = 5'b00000; w[173][34] = 5'b01111; w[173][35] = 5'b01111; w[173][36] = 5'b01111; w[173][37] = 5'b10000; w[173][38] = 5'b10000; w[173][39] = 5'b10000; w[173][40] = 5'b00000; w[173][41] = 5'b00000; w[173][42] = 5'b00000; w[173][43] = 5'b00000; w[173][44] = 5'b10000; w[173][45] = 5'b10000; w[173][46] = 5'b10000; w[173][47] = 5'b00000; w[173][48] = 5'b01111; w[173][49] = 5'b01111; w[173][50] = 5'b01111; w[173][51] = 5'b10000; w[173][52] = 5'b10000; w[173][53] = 5'b10000; w[173][54] = 5'b00000; w[173][55] = 5'b00000; w[173][56] = 5'b00000; w[173][57] = 5'b00000; w[173][58] = 5'b01111; w[173][59] = 5'b00000; w[173][60] = 5'b00000; w[173][61] = 5'b10000; w[173][62] = 5'b10000; w[173][63] = 5'b00000; w[173][64] = 5'b00000; w[173][65] = 5'b00000; w[173][66] = 5'b00000; w[173][67] = 5'b01111; w[173][68] = 5'b00000; w[173][69] = 5'b00000; w[173][70] = 5'b00000; w[173][71] = 5'b00000; w[173][72] = 5'b01111; w[173][73] = 5'b00000; w[173][74] = 5'b10000; w[173][75] = 5'b10000; w[173][76] = 5'b10000; w[173][77] = 5'b00000; w[173][78] = 5'b00000; w[173][79] = 5'b10000; w[173][80] = 5'b00000; w[173][81] = 5'b01111; w[173][82] = 5'b00000; w[173][83] = 5'b00000; w[173][84] = 5'b00000; w[173][85] = 5'b00000; w[173][86] = 5'b01111; w[173][87] = 5'b00000; w[173][88] = 5'b10000; w[173][89] = 5'b10000; w[173][90] = 5'b10000; w[173][91] = 5'b10000; w[173][92] = 5'b00000; w[173][93] = 5'b10000; w[173][94] = 5'b10000; w[173][95] = 5'b00000; w[173][96] = 5'b00000; w[173][97] = 5'b00000; w[173][98] = 5'b00000; w[173][99] = 5'b00000; w[173][100] = 5'b01111; w[173][101] = 5'b00000; w[173][102] = 5'b10000; w[173][103] = 5'b00000; w[173][104] = 5'b10000; w[173][105] = 5'b10000; w[173][106] = 5'b01111; w[173][107] = 5'b00000; w[173][108] = 5'b00000; w[173][109] = 5'b01111; w[173][110] = 5'b00000; w[173][111] = 5'b00000; w[173][112] = 5'b00000; w[173][113] = 5'b00000; w[173][114] = 5'b01111; w[173][115] = 5'b00000; w[173][116] = 5'b10000; w[173][117] = 5'b00000; w[173][118] = 5'b10000; w[173][119] = 5'b10000; w[173][120] = 5'b00000; w[173][121] = 5'b00000; w[173][122] = 5'b00000; w[173][123] = 5'b01111; w[173][124] = 5'b00000; w[173][125] = 5'b00000; w[173][126] = 5'b00000; w[173][127] = 5'b00000; w[173][128] = 5'b01111; w[173][129] = 5'b00000; w[173][130] = 5'b10000; w[173][131] = 5'b00000; w[173][132] = 5'b00000; w[173][133] = 5'b10000; w[173][134] = 5'b10000; w[173][135] = 5'b10000; w[173][136] = 5'b00000; w[173][137] = 5'b01111; w[173][138] = 5'b00000; w[173][139] = 5'b00000; w[173][140] = 5'b00000; w[173][141] = 5'b00000; w[173][142] = 5'b01111; w[173][143] = 5'b00000; w[173][144] = 5'b00000; w[173][145] = 5'b00000; w[173][146] = 5'b00000; w[173][147] = 5'b10000; w[173][148] = 5'b10000; w[173][149] = 5'b00000; w[173][150] = 5'b00000; w[173][151] = 5'b01111; w[173][152] = 5'b00000; w[173][153] = 5'b00000; w[173][154] = 5'b00000; w[173][155] = 5'b00000; w[173][156] = 5'b00000; w[173][157] = 5'b00000; w[173][158] = 5'b00000; w[173][159] = 5'b01111; w[173][160] = 5'b01111; w[173][161] = 5'b01111; w[173][162] = 5'b01111; w[173][163] = 5'b00000; w[173][164] = 5'b00000; w[173][165] = 5'b00000; w[173][166] = 5'b00000; w[173][167] = 5'b00000; w[173][168] = 5'b00000; w[173][169] = 5'b00000; w[173][170] = 5'b00000; w[173][171] = 5'b10000; w[173][172] = 5'b00000; w[173][173] = 5'b00000; w[173][174] = 5'b01111; w[173][175] = 5'b01111; w[173][176] = 5'b01111; w[173][177] = 5'b00000; w[173][178] = 5'b10000; w[173][179] = 5'b00000; w[173][180] = 5'b00000; w[173][181] = 5'b00000; w[173][182] = 5'b00000; w[173][183] = 5'b00000; w[173][184] = 5'b00000; w[173][185] = 5'b00000; w[173][186] = 5'b00000; w[173][187] = 5'b00000; w[173][188] = 5'b00000; w[173][189] = 5'b00000; w[173][190] = 5'b00000; w[173][191] = 5'b00000; w[173][192] = 5'b00000; w[173][193] = 5'b00000; w[173][194] = 5'b00000; w[173][195] = 5'b00000; w[173][196] = 5'b00000; w[173][197] = 5'b00000; w[173][198] = 5'b00000; w[173][199] = 5'b00000; w[173][200] = 5'b00000; w[173][201] = 5'b00000; w[173][202] = 5'b00000; w[173][203] = 5'b00000; w[173][204] = 5'b00000; w[173][205] = 5'b00000; w[173][206] = 5'b00000; w[173][207] = 5'b00000; w[173][208] = 5'b00000; w[173][209] = 5'b00000; 
w[174][0] = 5'b10000; w[174][1] = 5'b10000; w[174][2] = 5'b10000; w[174][3] = 5'b10000; w[174][4] = 5'b10000; w[174][5] = 5'b10000; w[174][6] = 5'b10000; w[174][7] = 5'b10000; w[174][8] = 5'b10000; w[174][9] = 5'b10000; w[174][10] = 5'b10000; w[174][11] = 5'b10000; w[174][12] = 5'b10000; w[174][13] = 5'b10000; w[174][14] = 5'b10000; w[174][15] = 5'b10000; w[174][16] = 5'b10000; w[174][17] = 5'b10000; w[174][18] = 5'b10000; w[174][19] = 5'b10000; w[174][20] = 5'b10000; w[174][21] = 5'b10000; w[174][22] = 5'b10000; w[174][23] = 5'b10000; w[174][24] = 5'b10000; w[174][25] = 5'b10000; w[174][26] = 5'b10000; w[174][27] = 5'b10000; w[174][28] = 5'b10000; w[174][29] = 5'b10000; w[174][30] = 5'b00000; w[174][31] = 5'b10000; w[174][32] = 5'b00000; w[174][33] = 5'b01111; w[174][34] = 5'b01111; w[174][35] = 5'b01111; w[174][36] = 5'b01111; w[174][37] = 5'b00000; w[174][38] = 5'b10000; w[174][39] = 5'b00000; w[174][40] = 5'b10000; w[174][41] = 5'b10000; w[174][42] = 5'b10000; w[174][43] = 5'b10000; w[174][44] = 5'b00000; w[174][45] = 5'b00000; w[174][46] = 5'b00000; w[174][47] = 5'b01111; w[174][48] = 5'b01111; w[174][49] = 5'b01111; w[174][50] = 5'b01111; w[174][51] = 5'b00000; w[174][52] = 5'b00000; w[174][53] = 5'b00000; w[174][54] = 5'b10000; w[174][55] = 5'b10000; w[174][56] = 5'b10000; w[174][57] = 5'b10000; w[174][58] = 5'b00000; w[174][59] = 5'b10000; w[174][60] = 5'b10000; w[174][61] = 5'b10000; w[174][62] = 5'b00000; w[174][63] = 5'b01111; w[174][64] = 5'b10000; w[174][65] = 5'b10000; w[174][66] = 5'b10000; w[174][67] = 5'b00000; w[174][68] = 5'b10000; w[174][69] = 5'b10000; w[174][70] = 5'b10000; w[174][71] = 5'b10000; w[174][72] = 5'b00000; w[174][73] = 5'b10000; w[174][74] = 5'b10000; w[174][75] = 5'b10000; w[174][76] = 5'b00000; w[174][77] = 5'b01111; w[174][78] = 5'b10000; w[174][79] = 5'b10000; w[174][80] = 5'b10000; w[174][81] = 5'b00000; w[174][82] = 5'b10000; w[174][83] = 5'b10000; w[174][84] = 5'b10000; w[174][85] = 5'b10000; w[174][86] = 5'b00000; w[174][87] = 5'b10000; w[174][88] = 5'b10000; w[174][89] = 5'b10000; w[174][90] = 5'b00000; w[174][91] = 5'b00000; w[174][92] = 5'b10000; w[174][93] = 5'b10000; w[174][94] = 5'b10000; w[174][95] = 5'b10000; w[174][96] = 5'b10000; w[174][97] = 5'b10000; w[174][98] = 5'b10000; w[174][99] = 5'b10000; w[174][100] = 5'b00000; w[174][101] = 5'b10000; w[174][102] = 5'b10000; w[174][103] = 5'b10000; w[174][104] = 5'b00000; w[174][105] = 5'b00000; w[174][106] = 5'b00000; w[174][107] = 5'b10000; w[174][108] = 5'b10000; w[174][109] = 5'b00000; w[174][110] = 5'b10000; w[174][111] = 5'b10000; w[174][112] = 5'b10000; w[174][113] = 5'b10000; w[174][114] = 5'b00000; w[174][115] = 5'b10000; w[174][116] = 5'b10000; w[174][117] = 5'b10000; w[174][118] = 5'b00000; w[174][119] = 5'b00000; w[174][120] = 5'b10000; w[174][121] = 5'b10000; w[174][122] = 5'b10000; w[174][123] = 5'b00000; w[174][124] = 5'b10000; w[174][125] = 5'b10000; w[174][126] = 5'b10000; w[174][127] = 5'b10000; w[174][128] = 5'b00000; w[174][129] = 5'b10000; w[174][130] = 5'b10000; w[174][131] = 5'b10000; w[174][132] = 5'b01111; w[174][133] = 5'b00000; w[174][134] = 5'b10000; w[174][135] = 5'b10000; w[174][136] = 5'b10000; w[174][137] = 5'b00000; w[174][138] = 5'b10000; w[174][139] = 5'b10000; w[174][140] = 5'b10000; w[174][141] = 5'b10000; w[174][142] = 5'b00000; w[174][143] = 5'b10000; w[174][144] = 5'b10000; w[174][145] = 5'b10000; w[174][146] = 5'b01111; w[174][147] = 5'b00000; w[174][148] = 5'b10000; w[174][149] = 5'b10000; w[174][150] = 5'b10000; w[174][151] = 5'b00000; w[174][152] = 5'b10000; w[174][153] = 5'b10000; w[174][154] = 5'b10000; w[174][155] = 5'b10000; w[174][156] = 5'b10000; w[174][157] = 5'b10000; w[174][158] = 5'b10000; w[174][159] = 5'b01111; w[174][160] = 5'b01111; w[174][161] = 5'b01111; w[174][162] = 5'b00000; w[174][163] = 5'b10000; w[174][164] = 5'b10000; w[174][165] = 5'b10000; w[174][166] = 5'b10000; w[174][167] = 5'b10000; w[174][168] = 5'b10000; w[174][169] = 5'b10000; w[174][170] = 5'b10000; w[174][171] = 5'b10000; w[174][172] = 5'b10000; w[174][173] = 5'b01111; w[174][174] = 5'b00000; w[174][175] = 5'b01111; w[174][176] = 5'b00000; w[174][177] = 5'b10000; w[174][178] = 5'b10000; w[174][179] = 5'b10000; w[174][180] = 5'b10000; w[174][181] = 5'b10000; w[174][182] = 5'b10000; w[174][183] = 5'b10000; w[174][184] = 5'b10000; w[174][185] = 5'b10000; w[174][186] = 5'b10000; w[174][187] = 5'b10000; w[174][188] = 5'b10000; w[174][189] = 5'b10000; w[174][190] = 5'b10000; w[174][191] = 5'b10000; w[174][192] = 5'b10000; w[174][193] = 5'b10000; w[174][194] = 5'b10000; w[174][195] = 5'b10000; w[174][196] = 5'b10000; w[174][197] = 5'b10000; w[174][198] = 5'b10000; w[174][199] = 5'b10000; w[174][200] = 5'b10000; w[174][201] = 5'b10000; w[174][202] = 5'b10000; w[174][203] = 5'b10000; w[174][204] = 5'b10000; w[174][205] = 5'b10000; w[174][206] = 5'b10000; w[174][207] = 5'b10000; w[174][208] = 5'b10000; w[174][209] = 5'b10000; 
w[175][0] = 5'b10000; w[175][1] = 5'b10000; w[175][2] = 5'b10000; w[175][3] = 5'b10000; w[175][4] = 5'b10000; w[175][5] = 5'b10000; w[175][6] = 5'b10000; w[175][7] = 5'b10000; w[175][8] = 5'b10000; w[175][9] = 5'b10000; w[175][10] = 5'b10000; w[175][11] = 5'b10000; w[175][12] = 5'b10000; w[175][13] = 5'b10000; w[175][14] = 5'b10000; w[175][15] = 5'b10000; w[175][16] = 5'b10000; w[175][17] = 5'b10000; w[175][18] = 5'b10000; w[175][19] = 5'b10000; w[175][20] = 5'b10000; w[175][21] = 5'b10000; w[175][22] = 5'b10000; w[175][23] = 5'b10000; w[175][24] = 5'b10000; w[175][25] = 5'b10000; w[175][26] = 5'b10000; w[175][27] = 5'b10000; w[175][28] = 5'b10000; w[175][29] = 5'b10000; w[175][30] = 5'b00000; w[175][31] = 5'b10000; w[175][32] = 5'b00000; w[175][33] = 5'b01111; w[175][34] = 5'b01111; w[175][35] = 5'b01111; w[175][36] = 5'b01111; w[175][37] = 5'b00000; w[175][38] = 5'b10000; w[175][39] = 5'b00000; w[175][40] = 5'b10000; w[175][41] = 5'b10000; w[175][42] = 5'b10000; w[175][43] = 5'b10000; w[175][44] = 5'b00000; w[175][45] = 5'b00000; w[175][46] = 5'b00000; w[175][47] = 5'b01111; w[175][48] = 5'b01111; w[175][49] = 5'b01111; w[175][50] = 5'b01111; w[175][51] = 5'b00000; w[175][52] = 5'b00000; w[175][53] = 5'b00000; w[175][54] = 5'b10000; w[175][55] = 5'b10000; w[175][56] = 5'b10000; w[175][57] = 5'b10000; w[175][58] = 5'b00000; w[175][59] = 5'b10000; w[175][60] = 5'b10000; w[175][61] = 5'b10000; w[175][62] = 5'b00000; w[175][63] = 5'b01111; w[175][64] = 5'b10000; w[175][65] = 5'b10000; w[175][66] = 5'b10000; w[175][67] = 5'b00000; w[175][68] = 5'b10000; w[175][69] = 5'b10000; w[175][70] = 5'b10000; w[175][71] = 5'b10000; w[175][72] = 5'b00000; w[175][73] = 5'b10000; w[175][74] = 5'b10000; w[175][75] = 5'b10000; w[175][76] = 5'b00000; w[175][77] = 5'b01111; w[175][78] = 5'b10000; w[175][79] = 5'b10000; w[175][80] = 5'b10000; w[175][81] = 5'b00000; w[175][82] = 5'b10000; w[175][83] = 5'b10000; w[175][84] = 5'b10000; w[175][85] = 5'b10000; w[175][86] = 5'b00000; w[175][87] = 5'b10000; w[175][88] = 5'b10000; w[175][89] = 5'b10000; w[175][90] = 5'b00000; w[175][91] = 5'b00000; w[175][92] = 5'b10000; w[175][93] = 5'b10000; w[175][94] = 5'b10000; w[175][95] = 5'b10000; w[175][96] = 5'b10000; w[175][97] = 5'b10000; w[175][98] = 5'b10000; w[175][99] = 5'b10000; w[175][100] = 5'b00000; w[175][101] = 5'b10000; w[175][102] = 5'b10000; w[175][103] = 5'b10000; w[175][104] = 5'b00000; w[175][105] = 5'b00000; w[175][106] = 5'b00000; w[175][107] = 5'b10000; w[175][108] = 5'b10000; w[175][109] = 5'b00000; w[175][110] = 5'b10000; w[175][111] = 5'b10000; w[175][112] = 5'b10000; w[175][113] = 5'b10000; w[175][114] = 5'b00000; w[175][115] = 5'b10000; w[175][116] = 5'b10000; w[175][117] = 5'b10000; w[175][118] = 5'b00000; w[175][119] = 5'b00000; w[175][120] = 5'b10000; w[175][121] = 5'b10000; w[175][122] = 5'b10000; w[175][123] = 5'b00000; w[175][124] = 5'b10000; w[175][125] = 5'b10000; w[175][126] = 5'b10000; w[175][127] = 5'b10000; w[175][128] = 5'b00000; w[175][129] = 5'b10000; w[175][130] = 5'b10000; w[175][131] = 5'b10000; w[175][132] = 5'b01111; w[175][133] = 5'b00000; w[175][134] = 5'b10000; w[175][135] = 5'b10000; w[175][136] = 5'b10000; w[175][137] = 5'b00000; w[175][138] = 5'b10000; w[175][139] = 5'b10000; w[175][140] = 5'b10000; w[175][141] = 5'b10000; w[175][142] = 5'b00000; w[175][143] = 5'b10000; w[175][144] = 5'b10000; w[175][145] = 5'b10000; w[175][146] = 5'b01111; w[175][147] = 5'b00000; w[175][148] = 5'b10000; w[175][149] = 5'b10000; w[175][150] = 5'b10000; w[175][151] = 5'b00000; w[175][152] = 5'b10000; w[175][153] = 5'b10000; w[175][154] = 5'b10000; w[175][155] = 5'b10000; w[175][156] = 5'b10000; w[175][157] = 5'b10000; w[175][158] = 5'b10000; w[175][159] = 5'b01111; w[175][160] = 5'b01111; w[175][161] = 5'b01111; w[175][162] = 5'b00000; w[175][163] = 5'b10000; w[175][164] = 5'b10000; w[175][165] = 5'b10000; w[175][166] = 5'b10000; w[175][167] = 5'b10000; w[175][168] = 5'b10000; w[175][169] = 5'b10000; w[175][170] = 5'b10000; w[175][171] = 5'b10000; w[175][172] = 5'b10000; w[175][173] = 5'b01111; w[175][174] = 5'b01111; w[175][175] = 5'b00000; w[175][176] = 5'b00000; w[175][177] = 5'b10000; w[175][178] = 5'b10000; w[175][179] = 5'b10000; w[175][180] = 5'b10000; w[175][181] = 5'b10000; w[175][182] = 5'b10000; w[175][183] = 5'b10000; w[175][184] = 5'b10000; w[175][185] = 5'b10000; w[175][186] = 5'b10000; w[175][187] = 5'b10000; w[175][188] = 5'b10000; w[175][189] = 5'b10000; w[175][190] = 5'b10000; w[175][191] = 5'b10000; w[175][192] = 5'b10000; w[175][193] = 5'b10000; w[175][194] = 5'b10000; w[175][195] = 5'b10000; w[175][196] = 5'b10000; w[175][197] = 5'b10000; w[175][198] = 5'b10000; w[175][199] = 5'b10000; w[175][200] = 5'b10000; w[175][201] = 5'b10000; w[175][202] = 5'b10000; w[175][203] = 5'b10000; w[175][204] = 5'b10000; w[175][205] = 5'b10000; w[175][206] = 5'b10000; w[175][207] = 5'b10000; w[175][208] = 5'b10000; w[175][209] = 5'b10000; 
w[176][0] = 5'b10000; w[176][1] = 5'b10000; w[176][2] = 5'b10000; w[176][3] = 5'b10000; w[176][4] = 5'b10000; w[176][5] = 5'b10000; w[176][6] = 5'b10000; w[176][7] = 5'b10000; w[176][8] = 5'b10000; w[176][9] = 5'b10000; w[176][10] = 5'b10000; w[176][11] = 5'b10000; w[176][12] = 5'b10000; w[176][13] = 5'b10000; w[176][14] = 5'b10000; w[176][15] = 5'b10000; w[176][16] = 5'b10000; w[176][17] = 5'b10000; w[176][18] = 5'b10000; w[176][19] = 5'b10000; w[176][20] = 5'b10000; w[176][21] = 5'b10000; w[176][22] = 5'b10000; w[176][23] = 5'b10000; w[176][24] = 5'b10000; w[176][25] = 5'b10000; w[176][26] = 5'b10000; w[176][27] = 5'b10000; w[176][28] = 5'b10000; w[176][29] = 5'b10000; w[176][30] = 5'b10000; w[176][31] = 5'b10000; w[176][32] = 5'b00000; w[176][33] = 5'b01111; w[176][34] = 5'b00000; w[176][35] = 5'b00000; w[176][36] = 5'b00000; w[176][37] = 5'b00000; w[176][38] = 5'b10000; w[176][39] = 5'b10000; w[176][40] = 5'b10000; w[176][41] = 5'b10000; w[176][42] = 5'b10000; w[176][43] = 5'b10000; w[176][44] = 5'b10000; w[176][45] = 5'b00000; w[176][46] = 5'b00000; w[176][47] = 5'b01111; w[176][48] = 5'b00000; w[176][49] = 5'b00000; w[176][50] = 5'b00000; w[176][51] = 5'b00000; w[176][52] = 5'b00000; w[176][53] = 5'b10000; w[176][54] = 5'b10000; w[176][55] = 5'b10000; w[176][56] = 5'b10000; w[176][57] = 5'b10000; w[176][58] = 5'b00000; w[176][59] = 5'b01111; w[176][60] = 5'b01111; w[176][61] = 5'b00000; w[176][62] = 5'b00000; w[176][63] = 5'b10000; w[176][64] = 5'b10000; w[176][65] = 5'b01111; w[176][66] = 5'b01111; w[176][67] = 5'b00000; w[176][68] = 5'b10000; w[176][69] = 5'b10000; w[176][70] = 5'b10000; w[176][71] = 5'b10000; w[176][72] = 5'b00000; w[176][73] = 5'b01111; w[176][74] = 5'b00000; w[176][75] = 5'b00000; w[176][76] = 5'b00000; w[176][77] = 5'b10000; w[176][78] = 5'b10000; w[176][79] = 5'b00000; w[176][80] = 5'b01111; w[176][81] = 5'b00000; w[176][82] = 5'b10000; w[176][83] = 5'b10000; w[176][84] = 5'b10000; w[176][85] = 5'b10000; w[176][86] = 5'b00000; w[176][87] = 5'b01111; w[176][88] = 5'b00000; w[176][89] = 5'b00000; w[176][90] = 5'b00000; w[176][91] = 5'b00000; w[176][92] = 5'b10000; w[176][93] = 5'b00000; w[176][94] = 5'b00000; w[176][95] = 5'b10000; w[176][96] = 5'b10000; w[176][97] = 5'b10000; w[176][98] = 5'b10000; w[176][99] = 5'b10000; w[176][100] = 5'b00000; w[176][101] = 5'b01111; w[176][102] = 5'b00000; w[176][103] = 5'b10000; w[176][104] = 5'b00000; w[176][105] = 5'b00000; w[176][106] = 5'b00000; w[176][107] = 5'b01111; w[176][108] = 5'b01111; w[176][109] = 5'b00000; w[176][110] = 5'b10000; w[176][111] = 5'b10000; w[176][112] = 5'b10000; w[176][113] = 5'b10000; w[176][114] = 5'b00000; w[176][115] = 5'b01111; w[176][116] = 5'b00000; w[176][117] = 5'b10000; w[176][118] = 5'b00000; w[176][119] = 5'b00000; w[176][120] = 5'b01111; w[176][121] = 5'b01111; w[176][122] = 5'b01111; w[176][123] = 5'b00000; w[176][124] = 5'b10000; w[176][125] = 5'b10000; w[176][126] = 5'b10000; w[176][127] = 5'b10000; w[176][128] = 5'b00000; w[176][129] = 5'b01111; w[176][130] = 5'b00000; w[176][131] = 5'b10000; w[176][132] = 5'b10000; w[176][133] = 5'b00000; w[176][134] = 5'b00000; w[176][135] = 5'b00000; w[176][136] = 5'b01111; w[176][137] = 5'b00000; w[176][138] = 5'b10000; w[176][139] = 5'b10000; w[176][140] = 5'b10000; w[176][141] = 5'b10000; w[176][142] = 5'b00000; w[176][143] = 5'b01111; w[176][144] = 5'b01111; w[176][145] = 5'b10000; w[176][146] = 5'b10000; w[176][147] = 5'b00000; w[176][148] = 5'b00000; w[176][149] = 5'b01111; w[176][150] = 5'b01111; w[176][151] = 5'b00000; w[176][152] = 5'b10000; w[176][153] = 5'b10000; w[176][154] = 5'b10000; w[176][155] = 5'b10000; w[176][156] = 5'b10000; w[176][157] = 5'b01111; w[176][158] = 5'b01111; w[176][159] = 5'b01111; w[176][160] = 5'b00000; w[176][161] = 5'b00000; w[176][162] = 5'b01111; w[176][163] = 5'b01111; w[176][164] = 5'b01111; w[176][165] = 5'b10000; w[176][166] = 5'b10000; w[176][167] = 5'b10000; w[176][168] = 5'b10000; w[176][169] = 5'b10000; w[176][170] = 5'b10000; w[176][171] = 5'b00000; w[176][172] = 5'b01111; w[176][173] = 5'b01111; w[176][174] = 5'b00000; w[176][175] = 5'b00000; w[176][176] = 5'b00000; w[176][177] = 5'b01111; w[176][178] = 5'b00000; w[176][179] = 5'b10000; w[176][180] = 5'b10000; w[176][181] = 5'b10000; w[176][182] = 5'b10000; w[176][183] = 5'b10000; w[176][184] = 5'b10000; w[176][185] = 5'b10000; w[176][186] = 5'b10000; w[176][187] = 5'b10000; w[176][188] = 5'b10000; w[176][189] = 5'b10000; w[176][190] = 5'b10000; w[176][191] = 5'b10000; w[176][192] = 5'b10000; w[176][193] = 5'b10000; w[176][194] = 5'b10000; w[176][195] = 5'b10000; w[176][196] = 5'b10000; w[176][197] = 5'b10000; w[176][198] = 5'b10000; w[176][199] = 5'b10000; w[176][200] = 5'b10000; w[176][201] = 5'b10000; w[176][202] = 5'b10000; w[176][203] = 5'b10000; w[176][204] = 5'b10000; w[176][205] = 5'b10000; w[176][206] = 5'b10000; w[176][207] = 5'b10000; w[176][208] = 5'b10000; w[176][209] = 5'b10000; 
w[177][0] = 5'b00000; w[177][1] = 5'b00000; w[177][2] = 5'b00000; w[177][3] = 5'b00000; w[177][4] = 5'b00000; w[177][5] = 5'b00000; w[177][6] = 5'b00000; w[177][7] = 5'b00000; w[177][8] = 5'b00000; w[177][9] = 5'b00000; w[177][10] = 5'b00000; w[177][11] = 5'b00000; w[177][12] = 5'b00000; w[177][13] = 5'b00000; w[177][14] = 5'b00000; w[177][15] = 5'b00000; w[177][16] = 5'b00000; w[177][17] = 5'b00000; w[177][18] = 5'b00000; w[177][19] = 5'b00000; w[177][20] = 5'b00000; w[177][21] = 5'b00000; w[177][22] = 5'b00000; w[177][23] = 5'b00000; w[177][24] = 5'b00000; w[177][25] = 5'b00000; w[177][26] = 5'b00000; w[177][27] = 5'b00000; w[177][28] = 5'b00000; w[177][29] = 5'b00000; w[177][30] = 5'b10000; w[177][31] = 5'b00000; w[177][32] = 5'b01111; w[177][33] = 5'b00000; w[177][34] = 5'b10000; w[177][35] = 5'b10000; w[177][36] = 5'b10000; w[177][37] = 5'b01111; w[177][38] = 5'b00000; w[177][39] = 5'b10000; w[177][40] = 5'b00000; w[177][41] = 5'b00000; w[177][42] = 5'b00000; w[177][43] = 5'b00000; w[177][44] = 5'b10000; w[177][45] = 5'b01111; w[177][46] = 5'b01111; w[177][47] = 5'b00000; w[177][48] = 5'b10000; w[177][49] = 5'b10000; w[177][50] = 5'b10000; w[177][51] = 5'b01111; w[177][52] = 5'b01111; w[177][53] = 5'b10000; w[177][54] = 5'b00000; w[177][55] = 5'b00000; w[177][56] = 5'b00000; w[177][57] = 5'b00000; w[177][58] = 5'b01111; w[177][59] = 5'b01111; w[177][60] = 5'b01111; w[177][61] = 5'b01111; w[177][62] = 5'b10000; w[177][63] = 5'b10000; w[177][64] = 5'b00000; w[177][65] = 5'b01111; w[177][66] = 5'b01111; w[177][67] = 5'b01111; w[177][68] = 5'b00000; w[177][69] = 5'b00000; w[177][70] = 5'b00000; w[177][71] = 5'b00000; w[177][72] = 5'b01111; w[177][73] = 5'b01111; w[177][74] = 5'b01111; w[177][75] = 5'b01111; w[177][76] = 5'b10000; w[177][77] = 5'b10000; w[177][78] = 5'b00000; w[177][79] = 5'b01111; w[177][80] = 5'b01111; w[177][81] = 5'b01111; w[177][82] = 5'b00000; w[177][83] = 5'b00000; w[177][84] = 5'b00000; w[177][85] = 5'b00000; w[177][86] = 5'b01111; w[177][87] = 5'b01111; w[177][88] = 5'b01111; w[177][89] = 5'b01111; w[177][90] = 5'b10000; w[177][91] = 5'b10000; w[177][92] = 5'b00000; w[177][93] = 5'b01111; w[177][94] = 5'b01111; w[177][95] = 5'b00000; w[177][96] = 5'b00000; w[177][97] = 5'b00000; w[177][98] = 5'b00000; w[177][99] = 5'b00000; w[177][100] = 5'b01111; w[177][101] = 5'b01111; w[177][102] = 5'b01111; w[177][103] = 5'b00000; w[177][104] = 5'b10000; w[177][105] = 5'b10000; w[177][106] = 5'b01111; w[177][107] = 5'b01111; w[177][108] = 5'b01111; w[177][109] = 5'b01111; w[177][110] = 5'b00000; w[177][111] = 5'b00000; w[177][112] = 5'b00000; w[177][113] = 5'b00000; w[177][114] = 5'b01111; w[177][115] = 5'b01111; w[177][116] = 5'b01111; w[177][117] = 5'b00000; w[177][118] = 5'b10000; w[177][119] = 5'b10000; w[177][120] = 5'b01111; w[177][121] = 5'b01111; w[177][122] = 5'b01111; w[177][123] = 5'b01111; w[177][124] = 5'b00000; w[177][125] = 5'b00000; w[177][126] = 5'b00000; w[177][127] = 5'b00000; w[177][128] = 5'b01111; w[177][129] = 5'b01111; w[177][130] = 5'b01111; w[177][131] = 5'b00000; w[177][132] = 5'b10000; w[177][133] = 5'b10000; w[177][134] = 5'b01111; w[177][135] = 5'b01111; w[177][136] = 5'b01111; w[177][137] = 5'b01111; w[177][138] = 5'b00000; w[177][139] = 5'b00000; w[177][140] = 5'b00000; w[177][141] = 5'b00000; w[177][142] = 5'b01111; w[177][143] = 5'b01111; w[177][144] = 5'b01111; w[177][145] = 5'b00000; w[177][146] = 5'b10000; w[177][147] = 5'b10000; w[177][148] = 5'b01111; w[177][149] = 5'b01111; w[177][150] = 5'b01111; w[177][151] = 5'b01111; w[177][152] = 5'b00000; w[177][153] = 5'b00000; w[177][154] = 5'b00000; w[177][155] = 5'b00000; w[177][156] = 5'b00000; w[177][157] = 5'b01111; w[177][158] = 5'b01111; w[177][159] = 5'b00000; w[177][160] = 5'b10000; w[177][161] = 5'b10000; w[177][162] = 5'b01111; w[177][163] = 5'b01111; w[177][164] = 5'b01111; w[177][165] = 5'b00000; w[177][166] = 5'b00000; w[177][167] = 5'b00000; w[177][168] = 5'b00000; w[177][169] = 5'b00000; w[177][170] = 5'b00000; w[177][171] = 5'b01111; w[177][172] = 5'b01111; w[177][173] = 5'b00000; w[177][174] = 5'b10000; w[177][175] = 5'b10000; w[177][176] = 5'b01111; w[177][177] = 5'b00000; w[177][178] = 5'b01111; w[177][179] = 5'b00000; w[177][180] = 5'b00000; w[177][181] = 5'b00000; w[177][182] = 5'b00000; w[177][183] = 5'b00000; w[177][184] = 5'b00000; w[177][185] = 5'b00000; w[177][186] = 5'b00000; w[177][187] = 5'b00000; w[177][188] = 5'b00000; w[177][189] = 5'b00000; w[177][190] = 5'b00000; w[177][191] = 5'b00000; w[177][192] = 5'b00000; w[177][193] = 5'b00000; w[177][194] = 5'b00000; w[177][195] = 5'b00000; w[177][196] = 5'b00000; w[177][197] = 5'b00000; w[177][198] = 5'b00000; w[177][199] = 5'b00000; w[177][200] = 5'b00000; w[177][201] = 5'b00000; w[177][202] = 5'b00000; w[177][203] = 5'b00000; w[177][204] = 5'b00000; w[177][205] = 5'b00000; w[177][206] = 5'b00000; w[177][207] = 5'b00000; w[177][208] = 5'b00000; w[177][209] = 5'b00000; 
w[178][0] = 5'b01111; w[178][1] = 5'b01111; w[178][2] = 5'b01111; w[178][3] = 5'b01111; w[178][4] = 5'b01111; w[178][5] = 5'b01111; w[178][6] = 5'b01111; w[178][7] = 5'b01111; w[178][8] = 5'b01111; w[178][9] = 5'b01111; w[178][10] = 5'b01111; w[178][11] = 5'b01111; w[178][12] = 5'b01111; w[178][13] = 5'b01111; w[178][14] = 5'b01111; w[178][15] = 5'b01111; w[178][16] = 5'b01111; w[178][17] = 5'b01111; w[178][18] = 5'b01111; w[178][19] = 5'b01111; w[178][20] = 5'b01111; w[178][21] = 5'b01111; w[178][22] = 5'b01111; w[178][23] = 5'b01111; w[178][24] = 5'b01111; w[178][25] = 5'b01111; w[178][26] = 5'b01111; w[178][27] = 5'b01111; w[178][28] = 5'b01111; w[178][29] = 5'b01111; w[178][30] = 5'b00000; w[178][31] = 5'b01111; w[178][32] = 5'b00000; w[178][33] = 5'b10000; w[178][34] = 5'b10000; w[178][35] = 5'b10000; w[178][36] = 5'b10000; w[178][37] = 5'b00000; w[178][38] = 5'b01111; w[178][39] = 5'b00000; w[178][40] = 5'b01111; w[178][41] = 5'b01111; w[178][42] = 5'b01111; w[178][43] = 5'b01111; w[178][44] = 5'b00000; w[178][45] = 5'b00000; w[178][46] = 5'b00000; w[178][47] = 5'b10000; w[178][48] = 5'b10000; w[178][49] = 5'b10000; w[178][50] = 5'b10000; w[178][51] = 5'b00000; w[178][52] = 5'b00000; w[178][53] = 5'b00000; w[178][54] = 5'b01111; w[178][55] = 5'b01111; w[178][56] = 5'b01111; w[178][57] = 5'b01111; w[178][58] = 5'b00000; w[178][59] = 5'b01111; w[178][60] = 5'b01111; w[178][61] = 5'b01111; w[178][62] = 5'b00000; w[178][63] = 5'b10000; w[178][64] = 5'b01111; w[178][65] = 5'b01111; w[178][66] = 5'b01111; w[178][67] = 5'b00000; w[178][68] = 5'b01111; w[178][69] = 5'b01111; w[178][70] = 5'b01111; w[178][71] = 5'b01111; w[178][72] = 5'b00000; w[178][73] = 5'b01111; w[178][74] = 5'b01111; w[178][75] = 5'b01111; w[178][76] = 5'b00000; w[178][77] = 5'b10000; w[178][78] = 5'b01111; w[178][79] = 5'b01111; w[178][80] = 5'b01111; w[178][81] = 5'b00000; w[178][82] = 5'b01111; w[178][83] = 5'b01111; w[178][84] = 5'b01111; w[178][85] = 5'b01111; w[178][86] = 5'b00000; w[178][87] = 5'b01111; w[178][88] = 5'b01111; w[178][89] = 5'b01111; w[178][90] = 5'b00000; w[178][91] = 5'b00000; w[178][92] = 5'b01111; w[178][93] = 5'b01111; w[178][94] = 5'b01111; w[178][95] = 5'b01111; w[178][96] = 5'b01111; w[178][97] = 5'b01111; w[178][98] = 5'b01111; w[178][99] = 5'b01111; w[178][100] = 5'b00000; w[178][101] = 5'b01111; w[178][102] = 5'b01111; w[178][103] = 5'b01111; w[178][104] = 5'b00000; w[178][105] = 5'b00000; w[178][106] = 5'b00000; w[178][107] = 5'b01111; w[178][108] = 5'b01111; w[178][109] = 5'b00000; w[178][110] = 5'b01111; w[178][111] = 5'b01111; w[178][112] = 5'b01111; w[178][113] = 5'b01111; w[178][114] = 5'b00000; w[178][115] = 5'b01111; w[178][116] = 5'b01111; w[178][117] = 5'b01111; w[178][118] = 5'b00000; w[178][119] = 5'b00000; w[178][120] = 5'b01111; w[178][121] = 5'b01111; w[178][122] = 5'b01111; w[178][123] = 5'b00000; w[178][124] = 5'b01111; w[178][125] = 5'b01111; w[178][126] = 5'b01111; w[178][127] = 5'b01111; w[178][128] = 5'b00000; w[178][129] = 5'b01111; w[178][130] = 5'b01111; w[178][131] = 5'b01111; w[178][132] = 5'b10000; w[178][133] = 5'b00000; w[178][134] = 5'b01111; w[178][135] = 5'b01111; w[178][136] = 5'b01111; w[178][137] = 5'b00000; w[178][138] = 5'b01111; w[178][139] = 5'b01111; w[178][140] = 5'b01111; w[178][141] = 5'b01111; w[178][142] = 5'b00000; w[178][143] = 5'b01111; w[178][144] = 5'b01111; w[178][145] = 5'b01111; w[178][146] = 5'b10000; w[178][147] = 5'b00000; w[178][148] = 5'b01111; w[178][149] = 5'b01111; w[178][150] = 5'b01111; w[178][151] = 5'b00000; w[178][152] = 5'b01111; w[178][153] = 5'b01111; w[178][154] = 5'b01111; w[178][155] = 5'b01111; w[178][156] = 5'b01111; w[178][157] = 5'b01111; w[178][158] = 5'b01111; w[178][159] = 5'b10000; w[178][160] = 5'b10000; w[178][161] = 5'b10000; w[178][162] = 5'b00000; w[178][163] = 5'b01111; w[178][164] = 5'b01111; w[178][165] = 5'b01111; w[178][166] = 5'b01111; w[178][167] = 5'b01111; w[178][168] = 5'b01111; w[178][169] = 5'b01111; w[178][170] = 5'b01111; w[178][171] = 5'b01111; w[178][172] = 5'b01111; w[178][173] = 5'b10000; w[178][174] = 5'b10000; w[178][175] = 5'b10000; w[178][176] = 5'b00000; w[178][177] = 5'b01111; w[178][178] = 5'b00000; w[178][179] = 5'b01111; w[178][180] = 5'b01111; w[178][181] = 5'b01111; w[178][182] = 5'b01111; w[178][183] = 5'b01111; w[178][184] = 5'b01111; w[178][185] = 5'b01111; w[178][186] = 5'b01111; w[178][187] = 5'b01111; w[178][188] = 5'b01111; w[178][189] = 5'b01111; w[178][190] = 5'b01111; w[178][191] = 5'b01111; w[178][192] = 5'b01111; w[178][193] = 5'b01111; w[178][194] = 5'b01111; w[178][195] = 5'b01111; w[178][196] = 5'b01111; w[178][197] = 5'b01111; w[178][198] = 5'b01111; w[178][199] = 5'b01111; w[178][200] = 5'b01111; w[178][201] = 5'b01111; w[178][202] = 5'b01111; w[178][203] = 5'b01111; w[178][204] = 5'b01111; w[178][205] = 5'b01111; w[178][206] = 5'b01111; w[178][207] = 5'b01111; w[178][208] = 5'b01111; w[178][209] = 5'b01111; 
w[179][0] = 5'b01111; w[179][1] = 5'b01111; w[179][2] = 5'b01111; w[179][3] = 5'b01111; w[179][4] = 5'b01111; w[179][5] = 5'b01111; w[179][6] = 5'b01111; w[179][7] = 5'b01111; w[179][8] = 5'b01111; w[179][9] = 5'b01111; w[179][10] = 5'b01111; w[179][11] = 5'b01111; w[179][12] = 5'b01111; w[179][13] = 5'b01111; w[179][14] = 5'b01111; w[179][15] = 5'b01111; w[179][16] = 5'b01111; w[179][17] = 5'b01111; w[179][18] = 5'b01111; w[179][19] = 5'b01111; w[179][20] = 5'b01111; w[179][21] = 5'b01111; w[179][22] = 5'b01111; w[179][23] = 5'b01111; w[179][24] = 5'b01111; w[179][25] = 5'b01111; w[179][26] = 5'b01111; w[179][27] = 5'b01111; w[179][28] = 5'b01111; w[179][29] = 5'b01111; w[179][30] = 5'b01111; w[179][31] = 5'b00000; w[179][32] = 5'b10000; w[179][33] = 5'b10000; w[179][34] = 5'b10000; w[179][35] = 5'b10000; w[179][36] = 5'b10000; w[179][37] = 5'b10000; w[179][38] = 5'b00000; w[179][39] = 5'b01111; w[179][40] = 5'b01111; w[179][41] = 5'b01111; w[179][42] = 5'b01111; w[179][43] = 5'b01111; w[179][44] = 5'b01111; w[179][45] = 5'b10000; w[179][46] = 5'b10000; w[179][47] = 5'b10000; w[179][48] = 5'b10000; w[179][49] = 5'b10000; w[179][50] = 5'b10000; w[179][51] = 5'b10000; w[179][52] = 5'b10000; w[179][53] = 5'b01111; w[179][54] = 5'b01111; w[179][55] = 5'b01111; w[179][56] = 5'b01111; w[179][57] = 5'b01111; w[179][58] = 5'b01111; w[179][59] = 5'b00000; w[179][60] = 5'b00000; w[179][61] = 5'b01111; w[179][62] = 5'b10000; w[179][63] = 5'b00000; w[179][64] = 5'b01111; w[179][65] = 5'b00000; w[179][66] = 5'b00000; w[179][67] = 5'b01111; w[179][68] = 5'b01111; w[179][69] = 5'b01111; w[179][70] = 5'b01111; w[179][71] = 5'b01111; w[179][72] = 5'b01111; w[179][73] = 5'b00000; w[179][74] = 5'b01111; w[179][75] = 5'b01111; w[179][76] = 5'b10000; w[179][77] = 5'b00000; w[179][78] = 5'b01111; w[179][79] = 5'b01111; w[179][80] = 5'b00000; w[179][81] = 5'b01111; w[179][82] = 5'b01111; w[179][83] = 5'b01111; w[179][84] = 5'b01111; w[179][85] = 5'b01111; w[179][86] = 5'b01111; w[179][87] = 5'b00000; w[179][88] = 5'b01111; w[179][89] = 5'b01111; w[179][90] = 5'b10000; w[179][91] = 5'b10000; w[179][92] = 5'b01111; w[179][93] = 5'b01111; w[179][94] = 5'b01111; w[179][95] = 5'b01111; w[179][96] = 5'b01111; w[179][97] = 5'b01111; w[179][98] = 5'b01111; w[179][99] = 5'b01111; w[179][100] = 5'b01111; w[179][101] = 5'b00000; w[179][102] = 5'b01111; w[179][103] = 5'b01111; w[179][104] = 5'b10000; w[179][105] = 5'b10000; w[179][106] = 5'b01111; w[179][107] = 5'b00000; w[179][108] = 5'b00000; w[179][109] = 5'b01111; w[179][110] = 5'b01111; w[179][111] = 5'b01111; w[179][112] = 5'b01111; w[179][113] = 5'b01111; w[179][114] = 5'b01111; w[179][115] = 5'b00000; w[179][116] = 5'b01111; w[179][117] = 5'b01111; w[179][118] = 5'b10000; w[179][119] = 5'b10000; w[179][120] = 5'b00000; w[179][121] = 5'b00000; w[179][122] = 5'b00000; w[179][123] = 5'b01111; w[179][124] = 5'b01111; w[179][125] = 5'b01111; w[179][126] = 5'b01111; w[179][127] = 5'b01111; w[179][128] = 5'b01111; w[179][129] = 5'b00000; w[179][130] = 5'b01111; w[179][131] = 5'b01111; w[179][132] = 5'b00000; w[179][133] = 5'b10000; w[179][134] = 5'b01111; w[179][135] = 5'b01111; w[179][136] = 5'b00000; w[179][137] = 5'b01111; w[179][138] = 5'b01111; w[179][139] = 5'b01111; w[179][140] = 5'b01111; w[179][141] = 5'b01111; w[179][142] = 5'b01111; w[179][143] = 5'b00000; w[179][144] = 5'b00000; w[179][145] = 5'b01111; w[179][146] = 5'b00000; w[179][147] = 5'b10000; w[179][148] = 5'b01111; w[179][149] = 5'b00000; w[179][150] = 5'b00000; w[179][151] = 5'b01111; w[179][152] = 5'b01111; w[179][153] = 5'b01111; w[179][154] = 5'b01111; w[179][155] = 5'b01111; w[179][156] = 5'b01111; w[179][157] = 5'b00000; w[179][158] = 5'b00000; w[179][159] = 5'b00000; w[179][160] = 5'b10000; w[179][161] = 5'b10000; w[179][162] = 5'b10000; w[179][163] = 5'b00000; w[179][164] = 5'b00000; w[179][165] = 5'b01111; w[179][166] = 5'b01111; w[179][167] = 5'b01111; w[179][168] = 5'b01111; w[179][169] = 5'b01111; w[179][170] = 5'b01111; w[179][171] = 5'b01111; w[179][172] = 5'b00000; w[179][173] = 5'b00000; w[179][174] = 5'b10000; w[179][175] = 5'b10000; w[179][176] = 5'b10000; w[179][177] = 5'b00000; w[179][178] = 5'b01111; w[179][179] = 5'b00000; w[179][180] = 5'b01111; w[179][181] = 5'b01111; w[179][182] = 5'b01111; w[179][183] = 5'b01111; w[179][184] = 5'b01111; w[179][185] = 5'b01111; w[179][186] = 5'b01111; w[179][187] = 5'b01111; w[179][188] = 5'b01111; w[179][189] = 5'b01111; w[179][190] = 5'b01111; w[179][191] = 5'b01111; w[179][192] = 5'b01111; w[179][193] = 5'b01111; w[179][194] = 5'b01111; w[179][195] = 5'b01111; w[179][196] = 5'b01111; w[179][197] = 5'b01111; w[179][198] = 5'b01111; w[179][199] = 5'b01111; w[179][200] = 5'b01111; w[179][201] = 5'b01111; w[179][202] = 5'b01111; w[179][203] = 5'b01111; w[179][204] = 5'b01111; w[179][205] = 5'b01111; w[179][206] = 5'b01111; w[179][207] = 5'b01111; w[179][208] = 5'b01111; w[179][209] = 5'b01111; 
w[180][0] = 5'b01111; w[180][1] = 5'b01111; w[180][2] = 5'b01111; w[180][3] = 5'b01111; w[180][4] = 5'b01111; w[180][5] = 5'b01111; w[180][6] = 5'b01111; w[180][7] = 5'b01111; w[180][8] = 5'b01111; w[180][9] = 5'b01111; w[180][10] = 5'b01111; w[180][11] = 5'b01111; w[180][12] = 5'b01111; w[180][13] = 5'b01111; w[180][14] = 5'b01111; w[180][15] = 5'b01111; w[180][16] = 5'b01111; w[180][17] = 5'b01111; w[180][18] = 5'b01111; w[180][19] = 5'b01111; w[180][20] = 5'b01111; w[180][21] = 5'b01111; w[180][22] = 5'b01111; w[180][23] = 5'b01111; w[180][24] = 5'b01111; w[180][25] = 5'b01111; w[180][26] = 5'b01111; w[180][27] = 5'b01111; w[180][28] = 5'b01111; w[180][29] = 5'b01111; w[180][30] = 5'b01111; w[180][31] = 5'b00000; w[180][32] = 5'b10000; w[180][33] = 5'b10000; w[180][34] = 5'b10000; w[180][35] = 5'b10000; w[180][36] = 5'b10000; w[180][37] = 5'b10000; w[180][38] = 5'b00000; w[180][39] = 5'b01111; w[180][40] = 5'b01111; w[180][41] = 5'b01111; w[180][42] = 5'b01111; w[180][43] = 5'b01111; w[180][44] = 5'b01111; w[180][45] = 5'b10000; w[180][46] = 5'b10000; w[180][47] = 5'b10000; w[180][48] = 5'b10000; w[180][49] = 5'b10000; w[180][50] = 5'b10000; w[180][51] = 5'b10000; w[180][52] = 5'b10000; w[180][53] = 5'b01111; w[180][54] = 5'b01111; w[180][55] = 5'b01111; w[180][56] = 5'b01111; w[180][57] = 5'b01111; w[180][58] = 5'b01111; w[180][59] = 5'b00000; w[180][60] = 5'b00000; w[180][61] = 5'b01111; w[180][62] = 5'b10000; w[180][63] = 5'b00000; w[180][64] = 5'b01111; w[180][65] = 5'b00000; w[180][66] = 5'b00000; w[180][67] = 5'b01111; w[180][68] = 5'b01111; w[180][69] = 5'b01111; w[180][70] = 5'b01111; w[180][71] = 5'b01111; w[180][72] = 5'b01111; w[180][73] = 5'b00000; w[180][74] = 5'b01111; w[180][75] = 5'b01111; w[180][76] = 5'b10000; w[180][77] = 5'b00000; w[180][78] = 5'b01111; w[180][79] = 5'b01111; w[180][80] = 5'b00000; w[180][81] = 5'b01111; w[180][82] = 5'b01111; w[180][83] = 5'b01111; w[180][84] = 5'b01111; w[180][85] = 5'b01111; w[180][86] = 5'b01111; w[180][87] = 5'b00000; w[180][88] = 5'b01111; w[180][89] = 5'b01111; w[180][90] = 5'b10000; w[180][91] = 5'b10000; w[180][92] = 5'b01111; w[180][93] = 5'b01111; w[180][94] = 5'b01111; w[180][95] = 5'b01111; w[180][96] = 5'b01111; w[180][97] = 5'b01111; w[180][98] = 5'b01111; w[180][99] = 5'b01111; w[180][100] = 5'b01111; w[180][101] = 5'b00000; w[180][102] = 5'b01111; w[180][103] = 5'b01111; w[180][104] = 5'b10000; w[180][105] = 5'b10000; w[180][106] = 5'b01111; w[180][107] = 5'b00000; w[180][108] = 5'b00000; w[180][109] = 5'b01111; w[180][110] = 5'b01111; w[180][111] = 5'b01111; w[180][112] = 5'b01111; w[180][113] = 5'b01111; w[180][114] = 5'b01111; w[180][115] = 5'b00000; w[180][116] = 5'b01111; w[180][117] = 5'b01111; w[180][118] = 5'b10000; w[180][119] = 5'b10000; w[180][120] = 5'b00000; w[180][121] = 5'b00000; w[180][122] = 5'b00000; w[180][123] = 5'b01111; w[180][124] = 5'b01111; w[180][125] = 5'b01111; w[180][126] = 5'b01111; w[180][127] = 5'b01111; w[180][128] = 5'b01111; w[180][129] = 5'b00000; w[180][130] = 5'b01111; w[180][131] = 5'b01111; w[180][132] = 5'b00000; w[180][133] = 5'b10000; w[180][134] = 5'b01111; w[180][135] = 5'b01111; w[180][136] = 5'b00000; w[180][137] = 5'b01111; w[180][138] = 5'b01111; w[180][139] = 5'b01111; w[180][140] = 5'b01111; w[180][141] = 5'b01111; w[180][142] = 5'b01111; w[180][143] = 5'b00000; w[180][144] = 5'b00000; w[180][145] = 5'b01111; w[180][146] = 5'b00000; w[180][147] = 5'b10000; w[180][148] = 5'b01111; w[180][149] = 5'b00000; w[180][150] = 5'b00000; w[180][151] = 5'b01111; w[180][152] = 5'b01111; w[180][153] = 5'b01111; w[180][154] = 5'b01111; w[180][155] = 5'b01111; w[180][156] = 5'b01111; w[180][157] = 5'b00000; w[180][158] = 5'b00000; w[180][159] = 5'b00000; w[180][160] = 5'b10000; w[180][161] = 5'b10000; w[180][162] = 5'b10000; w[180][163] = 5'b00000; w[180][164] = 5'b00000; w[180][165] = 5'b01111; w[180][166] = 5'b01111; w[180][167] = 5'b01111; w[180][168] = 5'b01111; w[180][169] = 5'b01111; w[180][170] = 5'b01111; w[180][171] = 5'b01111; w[180][172] = 5'b00000; w[180][173] = 5'b00000; w[180][174] = 5'b10000; w[180][175] = 5'b10000; w[180][176] = 5'b10000; w[180][177] = 5'b00000; w[180][178] = 5'b01111; w[180][179] = 5'b01111; w[180][180] = 5'b00000; w[180][181] = 5'b01111; w[180][182] = 5'b01111; w[180][183] = 5'b01111; w[180][184] = 5'b01111; w[180][185] = 5'b01111; w[180][186] = 5'b01111; w[180][187] = 5'b01111; w[180][188] = 5'b01111; w[180][189] = 5'b01111; w[180][190] = 5'b01111; w[180][191] = 5'b01111; w[180][192] = 5'b01111; w[180][193] = 5'b01111; w[180][194] = 5'b01111; w[180][195] = 5'b01111; w[180][196] = 5'b01111; w[180][197] = 5'b01111; w[180][198] = 5'b01111; w[180][199] = 5'b01111; w[180][200] = 5'b01111; w[180][201] = 5'b01111; w[180][202] = 5'b01111; w[180][203] = 5'b01111; w[180][204] = 5'b01111; w[180][205] = 5'b01111; w[180][206] = 5'b01111; w[180][207] = 5'b01111; w[180][208] = 5'b01111; w[180][209] = 5'b01111; 
w[181][0] = 5'b01111; w[181][1] = 5'b01111; w[181][2] = 5'b01111; w[181][3] = 5'b01111; w[181][4] = 5'b01111; w[181][5] = 5'b01111; w[181][6] = 5'b01111; w[181][7] = 5'b01111; w[181][8] = 5'b01111; w[181][9] = 5'b01111; w[181][10] = 5'b01111; w[181][11] = 5'b01111; w[181][12] = 5'b01111; w[181][13] = 5'b01111; w[181][14] = 5'b01111; w[181][15] = 5'b01111; w[181][16] = 5'b01111; w[181][17] = 5'b01111; w[181][18] = 5'b01111; w[181][19] = 5'b01111; w[181][20] = 5'b01111; w[181][21] = 5'b01111; w[181][22] = 5'b01111; w[181][23] = 5'b01111; w[181][24] = 5'b01111; w[181][25] = 5'b01111; w[181][26] = 5'b01111; w[181][27] = 5'b01111; w[181][28] = 5'b01111; w[181][29] = 5'b01111; w[181][30] = 5'b01111; w[181][31] = 5'b00000; w[181][32] = 5'b10000; w[181][33] = 5'b10000; w[181][34] = 5'b10000; w[181][35] = 5'b10000; w[181][36] = 5'b10000; w[181][37] = 5'b10000; w[181][38] = 5'b00000; w[181][39] = 5'b01111; w[181][40] = 5'b01111; w[181][41] = 5'b01111; w[181][42] = 5'b01111; w[181][43] = 5'b01111; w[181][44] = 5'b01111; w[181][45] = 5'b10000; w[181][46] = 5'b10000; w[181][47] = 5'b10000; w[181][48] = 5'b10000; w[181][49] = 5'b10000; w[181][50] = 5'b10000; w[181][51] = 5'b10000; w[181][52] = 5'b10000; w[181][53] = 5'b01111; w[181][54] = 5'b01111; w[181][55] = 5'b01111; w[181][56] = 5'b01111; w[181][57] = 5'b01111; w[181][58] = 5'b01111; w[181][59] = 5'b00000; w[181][60] = 5'b00000; w[181][61] = 5'b01111; w[181][62] = 5'b10000; w[181][63] = 5'b00000; w[181][64] = 5'b01111; w[181][65] = 5'b00000; w[181][66] = 5'b00000; w[181][67] = 5'b01111; w[181][68] = 5'b01111; w[181][69] = 5'b01111; w[181][70] = 5'b01111; w[181][71] = 5'b01111; w[181][72] = 5'b01111; w[181][73] = 5'b00000; w[181][74] = 5'b01111; w[181][75] = 5'b01111; w[181][76] = 5'b10000; w[181][77] = 5'b00000; w[181][78] = 5'b01111; w[181][79] = 5'b01111; w[181][80] = 5'b00000; w[181][81] = 5'b01111; w[181][82] = 5'b01111; w[181][83] = 5'b01111; w[181][84] = 5'b01111; w[181][85] = 5'b01111; w[181][86] = 5'b01111; w[181][87] = 5'b00000; w[181][88] = 5'b01111; w[181][89] = 5'b01111; w[181][90] = 5'b10000; w[181][91] = 5'b10000; w[181][92] = 5'b01111; w[181][93] = 5'b01111; w[181][94] = 5'b01111; w[181][95] = 5'b01111; w[181][96] = 5'b01111; w[181][97] = 5'b01111; w[181][98] = 5'b01111; w[181][99] = 5'b01111; w[181][100] = 5'b01111; w[181][101] = 5'b00000; w[181][102] = 5'b01111; w[181][103] = 5'b01111; w[181][104] = 5'b10000; w[181][105] = 5'b10000; w[181][106] = 5'b01111; w[181][107] = 5'b00000; w[181][108] = 5'b00000; w[181][109] = 5'b01111; w[181][110] = 5'b01111; w[181][111] = 5'b01111; w[181][112] = 5'b01111; w[181][113] = 5'b01111; w[181][114] = 5'b01111; w[181][115] = 5'b00000; w[181][116] = 5'b01111; w[181][117] = 5'b01111; w[181][118] = 5'b10000; w[181][119] = 5'b10000; w[181][120] = 5'b00000; w[181][121] = 5'b00000; w[181][122] = 5'b00000; w[181][123] = 5'b01111; w[181][124] = 5'b01111; w[181][125] = 5'b01111; w[181][126] = 5'b01111; w[181][127] = 5'b01111; w[181][128] = 5'b01111; w[181][129] = 5'b00000; w[181][130] = 5'b01111; w[181][131] = 5'b01111; w[181][132] = 5'b00000; w[181][133] = 5'b10000; w[181][134] = 5'b01111; w[181][135] = 5'b01111; w[181][136] = 5'b00000; w[181][137] = 5'b01111; w[181][138] = 5'b01111; w[181][139] = 5'b01111; w[181][140] = 5'b01111; w[181][141] = 5'b01111; w[181][142] = 5'b01111; w[181][143] = 5'b00000; w[181][144] = 5'b00000; w[181][145] = 5'b01111; w[181][146] = 5'b00000; w[181][147] = 5'b10000; w[181][148] = 5'b01111; w[181][149] = 5'b00000; w[181][150] = 5'b00000; w[181][151] = 5'b01111; w[181][152] = 5'b01111; w[181][153] = 5'b01111; w[181][154] = 5'b01111; w[181][155] = 5'b01111; w[181][156] = 5'b01111; w[181][157] = 5'b00000; w[181][158] = 5'b00000; w[181][159] = 5'b00000; w[181][160] = 5'b10000; w[181][161] = 5'b10000; w[181][162] = 5'b10000; w[181][163] = 5'b00000; w[181][164] = 5'b00000; w[181][165] = 5'b01111; w[181][166] = 5'b01111; w[181][167] = 5'b01111; w[181][168] = 5'b01111; w[181][169] = 5'b01111; w[181][170] = 5'b01111; w[181][171] = 5'b01111; w[181][172] = 5'b00000; w[181][173] = 5'b00000; w[181][174] = 5'b10000; w[181][175] = 5'b10000; w[181][176] = 5'b10000; w[181][177] = 5'b00000; w[181][178] = 5'b01111; w[181][179] = 5'b01111; w[181][180] = 5'b01111; w[181][181] = 5'b00000; w[181][182] = 5'b01111; w[181][183] = 5'b01111; w[181][184] = 5'b01111; w[181][185] = 5'b01111; w[181][186] = 5'b01111; w[181][187] = 5'b01111; w[181][188] = 5'b01111; w[181][189] = 5'b01111; w[181][190] = 5'b01111; w[181][191] = 5'b01111; w[181][192] = 5'b01111; w[181][193] = 5'b01111; w[181][194] = 5'b01111; w[181][195] = 5'b01111; w[181][196] = 5'b01111; w[181][197] = 5'b01111; w[181][198] = 5'b01111; w[181][199] = 5'b01111; w[181][200] = 5'b01111; w[181][201] = 5'b01111; w[181][202] = 5'b01111; w[181][203] = 5'b01111; w[181][204] = 5'b01111; w[181][205] = 5'b01111; w[181][206] = 5'b01111; w[181][207] = 5'b01111; w[181][208] = 5'b01111; w[181][209] = 5'b01111; 
w[182][0] = 5'b01111; w[182][1] = 5'b01111; w[182][2] = 5'b01111; w[182][3] = 5'b01111; w[182][4] = 5'b01111; w[182][5] = 5'b01111; w[182][6] = 5'b01111; w[182][7] = 5'b01111; w[182][8] = 5'b01111; w[182][9] = 5'b01111; w[182][10] = 5'b01111; w[182][11] = 5'b01111; w[182][12] = 5'b01111; w[182][13] = 5'b01111; w[182][14] = 5'b01111; w[182][15] = 5'b01111; w[182][16] = 5'b01111; w[182][17] = 5'b01111; w[182][18] = 5'b01111; w[182][19] = 5'b01111; w[182][20] = 5'b01111; w[182][21] = 5'b01111; w[182][22] = 5'b01111; w[182][23] = 5'b01111; w[182][24] = 5'b01111; w[182][25] = 5'b01111; w[182][26] = 5'b01111; w[182][27] = 5'b01111; w[182][28] = 5'b01111; w[182][29] = 5'b01111; w[182][30] = 5'b01111; w[182][31] = 5'b00000; w[182][32] = 5'b10000; w[182][33] = 5'b10000; w[182][34] = 5'b10000; w[182][35] = 5'b10000; w[182][36] = 5'b10000; w[182][37] = 5'b10000; w[182][38] = 5'b00000; w[182][39] = 5'b01111; w[182][40] = 5'b01111; w[182][41] = 5'b01111; w[182][42] = 5'b01111; w[182][43] = 5'b01111; w[182][44] = 5'b01111; w[182][45] = 5'b10000; w[182][46] = 5'b10000; w[182][47] = 5'b10000; w[182][48] = 5'b10000; w[182][49] = 5'b10000; w[182][50] = 5'b10000; w[182][51] = 5'b10000; w[182][52] = 5'b10000; w[182][53] = 5'b01111; w[182][54] = 5'b01111; w[182][55] = 5'b01111; w[182][56] = 5'b01111; w[182][57] = 5'b01111; w[182][58] = 5'b01111; w[182][59] = 5'b00000; w[182][60] = 5'b00000; w[182][61] = 5'b01111; w[182][62] = 5'b10000; w[182][63] = 5'b00000; w[182][64] = 5'b01111; w[182][65] = 5'b00000; w[182][66] = 5'b00000; w[182][67] = 5'b01111; w[182][68] = 5'b01111; w[182][69] = 5'b01111; w[182][70] = 5'b01111; w[182][71] = 5'b01111; w[182][72] = 5'b01111; w[182][73] = 5'b00000; w[182][74] = 5'b01111; w[182][75] = 5'b01111; w[182][76] = 5'b10000; w[182][77] = 5'b00000; w[182][78] = 5'b01111; w[182][79] = 5'b01111; w[182][80] = 5'b00000; w[182][81] = 5'b01111; w[182][82] = 5'b01111; w[182][83] = 5'b01111; w[182][84] = 5'b01111; w[182][85] = 5'b01111; w[182][86] = 5'b01111; w[182][87] = 5'b00000; w[182][88] = 5'b01111; w[182][89] = 5'b01111; w[182][90] = 5'b10000; w[182][91] = 5'b10000; w[182][92] = 5'b01111; w[182][93] = 5'b01111; w[182][94] = 5'b01111; w[182][95] = 5'b01111; w[182][96] = 5'b01111; w[182][97] = 5'b01111; w[182][98] = 5'b01111; w[182][99] = 5'b01111; w[182][100] = 5'b01111; w[182][101] = 5'b00000; w[182][102] = 5'b01111; w[182][103] = 5'b01111; w[182][104] = 5'b10000; w[182][105] = 5'b10000; w[182][106] = 5'b01111; w[182][107] = 5'b00000; w[182][108] = 5'b00000; w[182][109] = 5'b01111; w[182][110] = 5'b01111; w[182][111] = 5'b01111; w[182][112] = 5'b01111; w[182][113] = 5'b01111; w[182][114] = 5'b01111; w[182][115] = 5'b00000; w[182][116] = 5'b01111; w[182][117] = 5'b01111; w[182][118] = 5'b10000; w[182][119] = 5'b10000; w[182][120] = 5'b00000; w[182][121] = 5'b00000; w[182][122] = 5'b00000; w[182][123] = 5'b01111; w[182][124] = 5'b01111; w[182][125] = 5'b01111; w[182][126] = 5'b01111; w[182][127] = 5'b01111; w[182][128] = 5'b01111; w[182][129] = 5'b00000; w[182][130] = 5'b01111; w[182][131] = 5'b01111; w[182][132] = 5'b00000; w[182][133] = 5'b10000; w[182][134] = 5'b01111; w[182][135] = 5'b01111; w[182][136] = 5'b00000; w[182][137] = 5'b01111; w[182][138] = 5'b01111; w[182][139] = 5'b01111; w[182][140] = 5'b01111; w[182][141] = 5'b01111; w[182][142] = 5'b01111; w[182][143] = 5'b00000; w[182][144] = 5'b00000; w[182][145] = 5'b01111; w[182][146] = 5'b00000; w[182][147] = 5'b10000; w[182][148] = 5'b01111; w[182][149] = 5'b00000; w[182][150] = 5'b00000; w[182][151] = 5'b01111; w[182][152] = 5'b01111; w[182][153] = 5'b01111; w[182][154] = 5'b01111; w[182][155] = 5'b01111; w[182][156] = 5'b01111; w[182][157] = 5'b00000; w[182][158] = 5'b00000; w[182][159] = 5'b00000; w[182][160] = 5'b10000; w[182][161] = 5'b10000; w[182][162] = 5'b10000; w[182][163] = 5'b00000; w[182][164] = 5'b00000; w[182][165] = 5'b01111; w[182][166] = 5'b01111; w[182][167] = 5'b01111; w[182][168] = 5'b01111; w[182][169] = 5'b01111; w[182][170] = 5'b01111; w[182][171] = 5'b01111; w[182][172] = 5'b00000; w[182][173] = 5'b00000; w[182][174] = 5'b10000; w[182][175] = 5'b10000; w[182][176] = 5'b10000; w[182][177] = 5'b00000; w[182][178] = 5'b01111; w[182][179] = 5'b01111; w[182][180] = 5'b01111; w[182][181] = 5'b01111; w[182][182] = 5'b00000; w[182][183] = 5'b01111; w[182][184] = 5'b01111; w[182][185] = 5'b01111; w[182][186] = 5'b01111; w[182][187] = 5'b01111; w[182][188] = 5'b01111; w[182][189] = 5'b01111; w[182][190] = 5'b01111; w[182][191] = 5'b01111; w[182][192] = 5'b01111; w[182][193] = 5'b01111; w[182][194] = 5'b01111; w[182][195] = 5'b01111; w[182][196] = 5'b01111; w[182][197] = 5'b01111; w[182][198] = 5'b01111; w[182][199] = 5'b01111; w[182][200] = 5'b01111; w[182][201] = 5'b01111; w[182][202] = 5'b01111; w[182][203] = 5'b01111; w[182][204] = 5'b01111; w[182][205] = 5'b01111; w[182][206] = 5'b01111; w[182][207] = 5'b01111; w[182][208] = 5'b01111; w[182][209] = 5'b01111; 
w[183][0] = 5'b01111; w[183][1] = 5'b01111; w[183][2] = 5'b01111; w[183][3] = 5'b01111; w[183][4] = 5'b01111; w[183][5] = 5'b01111; w[183][6] = 5'b01111; w[183][7] = 5'b01111; w[183][8] = 5'b01111; w[183][9] = 5'b01111; w[183][10] = 5'b01111; w[183][11] = 5'b01111; w[183][12] = 5'b01111; w[183][13] = 5'b01111; w[183][14] = 5'b01111; w[183][15] = 5'b01111; w[183][16] = 5'b01111; w[183][17] = 5'b01111; w[183][18] = 5'b01111; w[183][19] = 5'b01111; w[183][20] = 5'b01111; w[183][21] = 5'b01111; w[183][22] = 5'b01111; w[183][23] = 5'b01111; w[183][24] = 5'b01111; w[183][25] = 5'b01111; w[183][26] = 5'b01111; w[183][27] = 5'b01111; w[183][28] = 5'b01111; w[183][29] = 5'b01111; w[183][30] = 5'b01111; w[183][31] = 5'b00000; w[183][32] = 5'b10000; w[183][33] = 5'b10000; w[183][34] = 5'b10000; w[183][35] = 5'b10000; w[183][36] = 5'b10000; w[183][37] = 5'b10000; w[183][38] = 5'b00000; w[183][39] = 5'b01111; w[183][40] = 5'b01111; w[183][41] = 5'b01111; w[183][42] = 5'b01111; w[183][43] = 5'b01111; w[183][44] = 5'b01111; w[183][45] = 5'b10000; w[183][46] = 5'b10000; w[183][47] = 5'b10000; w[183][48] = 5'b10000; w[183][49] = 5'b10000; w[183][50] = 5'b10000; w[183][51] = 5'b10000; w[183][52] = 5'b10000; w[183][53] = 5'b01111; w[183][54] = 5'b01111; w[183][55] = 5'b01111; w[183][56] = 5'b01111; w[183][57] = 5'b01111; w[183][58] = 5'b01111; w[183][59] = 5'b00000; w[183][60] = 5'b00000; w[183][61] = 5'b01111; w[183][62] = 5'b10000; w[183][63] = 5'b00000; w[183][64] = 5'b01111; w[183][65] = 5'b00000; w[183][66] = 5'b00000; w[183][67] = 5'b01111; w[183][68] = 5'b01111; w[183][69] = 5'b01111; w[183][70] = 5'b01111; w[183][71] = 5'b01111; w[183][72] = 5'b01111; w[183][73] = 5'b00000; w[183][74] = 5'b01111; w[183][75] = 5'b01111; w[183][76] = 5'b10000; w[183][77] = 5'b00000; w[183][78] = 5'b01111; w[183][79] = 5'b01111; w[183][80] = 5'b00000; w[183][81] = 5'b01111; w[183][82] = 5'b01111; w[183][83] = 5'b01111; w[183][84] = 5'b01111; w[183][85] = 5'b01111; w[183][86] = 5'b01111; w[183][87] = 5'b00000; w[183][88] = 5'b01111; w[183][89] = 5'b01111; w[183][90] = 5'b10000; w[183][91] = 5'b10000; w[183][92] = 5'b01111; w[183][93] = 5'b01111; w[183][94] = 5'b01111; w[183][95] = 5'b01111; w[183][96] = 5'b01111; w[183][97] = 5'b01111; w[183][98] = 5'b01111; w[183][99] = 5'b01111; w[183][100] = 5'b01111; w[183][101] = 5'b00000; w[183][102] = 5'b01111; w[183][103] = 5'b01111; w[183][104] = 5'b10000; w[183][105] = 5'b10000; w[183][106] = 5'b01111; w[183][107] = 5'b00000; w[183][108] = 5'b00000; w[183][109] = 5'b01111; w[183][110] = 5'b01111; w[183][111] = 5'b01111; w[183][112] = 5'b01111; w[183][113] = 5'b01111; w[183][114] = 5'b01111; w[183][115] = 5'b00000; w[183][116] = 5'b01111; w[183][117] = 5'b01111; w[183][118] = 5'b10000; w[183][119] = 5'b10000; w[183][120] = 5'b00000; w[183][121] = 5'b00000; w[183][122] = 5'b00000; w[183][123] = 5'b01111; w[183][124] = 5'b01111; w[183][125] = 5'b01111; w[183][126] = 5'b01111; w[183][127] = 5'b01111; w[183][128] = 5'b01111; w[183][129] = 5'b00000; w[183][130] = 5'b01111; w[183][131] = 5'b01111; w[183][132] = 5'b00000; w[183][133] = 5'b10000; w[183][134] = 5'b01111; w[183][135] = 5'b01111; w[183][136] = 5'b00000; w[183][137] = 5'b01111; w[183][138] = 5'b01111; w[183][139] = 5'b01111; w[183][140] = 5'b01111; w[183][141] = 5'b01111; w[183][142] = 5'b01111; w[183][143] = 5'b00000; w[183][144] = 5'b00000; w[183][145] = 5'b01111; w[183][146] = 5'b00000; w[183][147] = 5'b10000; w[183][148] = 5'b01111; w[183][149] = 5'b00000; w[183][150] = 5'b00000; w[183][151] = 5'b01111; w[183][152] = 5'b01111; w[183][153] = 5'b01111; w[183][154] = 5'b01111; w[183][155] = 5'b01111; w[183][156] = 5'b01111; w[183][157] = 5'b00000; w[183][158] = 5'b00000; w[183][159] = 5'b00000; w[183][160] = 5'b10000; w[183][161] = 5'b10000; w[183][162] = 5'b10000; w[183][163] = 5'b00000; w[183][164] = 5'b00000; w[183][165] = 5'b01111; w[183][166] = 5'b01111; w[183][167] = 5'b01111; w[183][168] = 5'b01111; w[183][169] = 5'b01111; w[183][170] = 5'b01111; w[183][171] = 5'b01111; w[183][172] = 5'b00000; w[183][173] = 5'b00000; w[183][174] = 5'b10000; w[183][175] = 5'b10000; w[183][176] = 5'b10000; w[183][177] = 5'b00000; w[183][178] = 5'b01111; w[183][179] = 5'b01111; w[183][180] = 5'b01111; w[183][181] = 5'b01111; w[183][182] = 5'b01111; w[183][183] = 5'b00000; w[183][184] = 5'b01111; w[183][185] = 5'b01111; w[183][186] = 5'b01111; w[183][187] = 5'b01111; w[183][188] = 5'b01111; w[183][189] = 5'b01111; w[183][190] = 5'b01111; w[183][191] = 5'b01111; w[183][192] = 5'b01111; w[183][193] = 5'b01111; w[183][194] = 5'b01111; w[183][195] = 5'b01111; w[183][196] = 5'b01111; w[183][197] = 5'b01111; w[183][198] = 5'b01111; w[183][199] = 5'b01111; w[183][200] = 5'b01111; w[183][201] = 5'b01111; w[183][202] = 5'b01111; w[183][203] = 5'b01111; w[183][204] = 5'b01111; w[183][205] = 5'b01111; w[183][206] = 5'b01111; w[183][207] = 5'b01111; w[183][208] = 5'b01111; w[183][209] = 5'b01111; 
w[184][0] = 5'b01111; w[184][1] = 5'b01111; w[184][2] = 5'b01111; w[184][3] = 5'b01111; w[184][4] = 5'b01111; w[184][5] = 5'b01111; w[184][6] = 5'b01111; w[184][7] = 5'b01111; w[184][8] = 5'b01111; w[184][9] = 5'b01111; w[184][10] = 5'b01111; w[184][11] = 5'b01111; w[184][12] = 5'b01111; w[184][13] = 5'b01111; w[184][14] = 5'b01111; w[184][15] = 5'b01111; w[184][16] = 5'b01111; w[184][17] = 5'b01111; w[184][18] = 5'b01111; w[184][19] = 5'b01111; w[184][20] = 5'b01111; w[184][21] = 5'b01111; w[184][22] = 5'b01111; w[184][23] = 5'b01111; w[184][24] = 5'b01111; w[184][25] = 5'b01111; w[184][26] = 5'b01111; w[184][27] = 5'b01111; w[184][28] = 5'b01111; w[184][29] = 5'b01111; w[184][30] = 5'b01111; w[184][31] = 5'b00000; w[184][32] = 5'b10000; w[184][33] = 5'b10000; w[184][34] = 5'b10000; w[184][35] = 5'b10000; w[184][36] = 5'b10000; w[184][37] = 5'b10000; w[184][38] = 5'b00000; w[184][39] = 5'b01111; w[184][40] = 5'b01111; w[184][41] = 5'b01111; w[184][42] = 5'b01111; w[184][43] = 5'b01111; w[184][44] = 5'b01111; w[184][45] = 5'b10000; w[184][46] = 5'b10000; w[184][47] = 5'b10000; w[184][48] = 5'b10000; w[184][49] = 5'b10000; w[184][50] = 5'b10000; w[184][51] = 5'b10000; w[184][52] = 5'b10000; w[184][53] = 5'b01111; w[184][54] = 5'b01111; w[184][55] = 5'b01111; w[184][56] = 5'b01111; w[184][57] = 5'b01111; w[184][58] = 5'b01111; w[184][59] = 5'b00000; w[184][60] = 5'b00000; w[184][61] = 5'b01111; w[184][62] = 5'b10000; w[184][63] = 5'b00000; w[184][64] = 5'b01111; w[184][65] = 5'b00000; w[184][66] = 5'b00000; w[184][67] = 5'b01111; w[184][68] = 5'b01111; w[184][69] = 5'b01111; w[184][70] = 5'b01111; w[184][71] = 5'b01111; w[184][72] = 5'b01111; w[184][73] = 5'b00000; w[184][74] = 5'b01111; w[184][75] = 5'b01111; w[184][76] = 5'b10000; w[184][77] = 5'b00000; w[184][78] = 5'b01111; w[184][79] = 5'b01111; w[184][80] = 5'b00000; w[184][81] = 5'b01111; w[184][82] = 5'b01111; w[184][83] = 5'b01111; w[184][84] = 5'b01111; w[184][85] = 5'b01111; w[184][86] = 5'b01111; w[184][87] = 5'b00000; w[184][88] = 5'b01111; w[184][89] = 5'b01111; w[184][90] = 5'b10000; w[184][91] = 5'b10000; w[184][92] = 5'b01111; w[184][93] = 5'b01111; w[184][94] = 5'b01111; w[184][95] = 5'b01111; w[184][96] = 5'b01111; w[184][97] = 5'b01111; w[184][98] = 5'b01111; w[184][99] = 5'b01111; w[184][100] = 5'b01111; w[184][101] = 5'b00000; w[184][102] = 5'b01111; w[184][103] = 5'b01111; w[184][104] = 5'b10000; w[184][105] = 5'b10000; w[184][106] = 5'b01111; w[184][107] = 5'b00000; w[184][108] = 5'b00000; w[184][109] = 5'b01111; w[184][110] = 5'b01111; w[184][111] = 5'b01111; w[184][112] = 5'b01111; w[184][113] = 5'b01111; w[184][114] = 5'b01111; w[184][115] = 5'b00000; w[184][116] = 5'b01111; w[184][117] = 5'b01111; w[184][118] = 5'b10000; w[184][119] = 5'b10000; w[184][120] = 5'b00000; w[184][121] = 5'b00000; w[184][122] = 5'b00000; w[184][123] = 5'b01111; w[184][124] = 5'b01111; w[184][125] = 5'b01111; w[184][126] = 5'b01111; w[184][127] = 5'b01111; w[184][128] = 5'b01111; w[184][129] = 5'b00000; w[184][130] = 5'b01111; w[184][131] = 5'b01111; w[184][132] = 5'b00000; w[184][133] = 5'b10000; w[184][134] = 5'b01111; w[184][135] = 5'b01111; w[184][136] = 5'b00000; w[184][137] = 5'b01111; w[184][138] = 5'b01111; w[184][139] = 5'b01111; w[184][140] = 5'b01111; w[184][141] = 5'b01111; w[184][142] = 5'b01111; w[184][143] = 5'b00000; w[184][144] = 5'b00000; w[184][145] = 5'b01111; w[184][146] = 5'b00000; w[184][147] = 5'b10000; w[184][148] = 5'b01111; w[184][149] = 5'b00000; w[184][150] = 5'b00000; w[184][151] = 5'b01111; w[184][152] = 5'b01111; w[184][153] = 5'b01111; w[184][154] = 5'b01111; w[184][155] = 5'b01111; w[184][156] = 5'b01111; w[184][157] = 5'b00000; w[184][158] = 5'b00000; w[184][159] = 5'b00000; w[184][160] = 5'b10000; w[184][161] = 5'b10000; w[184][162] = 5'b10000; w[184][163] = 5'b00000; w[184][164] = 5'b00000; w[184][165] = 5'b01111; w[184][166] = 5'b01111; w[184][167] = 5'b01111; w[184][168] = 5'b01111; w[184][169] = 5'b01111; w[184][170] = 5'b01111; w[184][171] = 5'b01111; w[184][172] = 5'b00000; w[184][173] = 5'b00000; w[184][174] = 5'b10000; w[184][175] = 5'b10000; w[184][176] = 5'b10000; w[184][177] = 5'b00000; w[184][178] = 5'b01111; w[184][179] = 5'b01111; w[184][180] = 5'b01111; w[184][181] = 5'b01111; w[184][182] = 5'b01111; w[184][183] = 5'b01111; w[184][184] = 5'b00000; w[184][185] = 5'b01111; w[184][186] = 5'b01111; w[184][187] = 5'b01111; w[184][188] = 5'b01111; w[184][189] = 5'b01111; w[184][190] = 5'b01111; w[184][191] = 5'b01111; w[184][192] = 5'b01111; w[184][193] = 5'b01111; w[184][194] = 5'b01111; w[184][195] = 5'b01111; w[184][196] = 5'b01111; w[184][197] = 5'b01111; w[184][198] = 5'b01111; w[184][199] = 5'b01111; w[184][200] = 5'b01111; w[184][201] = 5'b01111; w[184][202] = 5'b01111; w[184][203] = 5'b01111; w[184][204] = 5'b01111; w[184][205] = 5'b01111; w[184][206] = 5'b01111; w[184][207] = 5'b01111; w[184][208] = 5'b01111; w[184][209] = 5'b01111; 
w[185][0] = 5'b01111; w[185][1] = 5'b01111; w[185][2] = 5'b01111; w[185][3] = 5'b01111; w[185][4] = 5'b01111; w[185][5] = 5'b01111; w[185][6] = 5'b01111; w[185][7] = 5'b01111; w[185][8] = 5'b01111; w[185][9] = 5'b01111; w[185][10] = 5'b01111; w[185][11] = 5'b01111; w[185][12] = 5'b01111; w[185][13] = 5'b01111; w[185][14] = 5'b01111; w[185][15] = 5'b01111; w[185][16] = 5'b01111; w[185][17] = 5'b01111; w[185][18] = 5'b01111; w[185][19] = 5'b01111; w[185][20] = 5'b01111; w[185][21] = 5'b01111; w[185][22] = 5'b01111; w[185][23] = 5'b01111; w[185][24] = 5'b01111; w[185][25] = 5'b01111; w[185][26] = 5'b01111; w[185][27] = 5'b01111; w[185][28] = 5'b01111; w[185][29] = 5'b01111; w[185][30] = 5'b01111; w[185][31] = 5'b00000; w[185][32] = 5'b10000; w[185][33] = 5'b10000; w[185][34] = 5'b10000; w[185][35] = 5'b10000; w[185][36] = 5'b10000; w[185][37] = 5'b10000; w[185][38] = 5'b00000; w[185][39] = 5'b01111; w[185][40] = 5'b01111; w[185][41] = 5'b01111; w[185][42] = 5'b01111; w[185][43] = 5'b01111; w[185][44] = 5'b01111; w[185][45] = 5'b10000; w[185][46] = 5'b10000; w[185][47] = 5'b10000; w[185][48] = 5'b10000; w[185][49] = 5'b10000; w[185][50] = 5'b10000; w[185][51] = 5'b10000; w[185][52] = 5'b10000; w[185][53] = 5'b01111; w[185][54] = 5'b01111; w[185][55] = 5'b01111; w[185][56] = 5'b01111; w[185][57] = 5'b01111; w[185][58] = 5'b01111; w[185][59] = 5'b00000; w[185][60] = 5'b00000; w[185][61] = 5'b01111; w[185][62] = 5'b10000; w[185][63] = 5'b00000; w[185][64] = 5'b01111; w[185][65] = 5'b00000; w[185][66] = 5'b00000; w[185][67] = 5'b01111; w[185][68] = 5'b01111; w[185][69] = 5'b01111; w[185][70] = 5'b01111; w[185][71] = 5'b01111; w[185][72] = 5'b01111; w[185][73] = 5'b00000; w[185][74] = 5'b01111; w[185][75] = 5'b01111; w[185][76] = 5'b10000; w[185][77] = 5'b00000; w[185][78] = 5'b01111; w[185][79] = 5'b01111; w[185][80] = 5'b00000; w[185][81] = 5'b01111; w[185][82] = 5'b01111; w[185][83] = 5'b01111; w[185][84] = 5'b01111; w[185][85] = 5'b01111; w[185][86] = 5'b01111; w[185][87] = 5'b00000; w[185][88] = 5'b01111; w[185][89] = 5'b01111; w[185][90] = 5'b10000; w[185][91] = 5'b10000; w[185][92] = 5'b01111; w[185][93] = 5'b01111; w[185][94] = 5'b01111; w[185][95] = 5'b01111; w[185][96] = 5'b01111; w[185][97] = 5'b01111; w[185][98] = 5'b01111; w[185][99] = 5'b01111; w[185][100] = 5'b01111; w[185][101] = 5'b00000; w[185][102] = 5'b01111; w[185][103] = 5'b01111; w[185][104] = 5'b10000; w[185][105] = 5'b10000; w[185][106] = 5'b01111; w[185][107] = 5'b00000; w[185][108] = 5'b00000; w[185][109] = 5'b01111; w[185][110] = 5'b01111; w[185][111] = 5'b01111; w[185][112] = 5'b01111; w[185][113] = 5'b01111; w[185][114] = 5'b01111; w[185][115] = 5'b00000; w[185][116] = 5'b01111; w[185][117] = 5'b01111; w[185][118] = 5'b10000; w[185][119] = 5'b10000; w[185][120] = 5'b00000; w[185][121] = 5'b00000; w[185][122] = 5'b00000; w[185][123] = 5'b01111; w[185][124] = 5'b01111; w[185][125] = 5'b01111; w[185][126] = 5'b01111; w[185][127] = 5'b01111; w[185][128] = 5'b01111; w[185][129] = 5'b00000; w[185][130] = 5'b01111; w[185][131] = 5'b01111; w[185][132] = 5'b00000; w[185][133] = 5'b10000; w[185][134] = 5'b01111; w[185][135] = 5'b01111; w[185][136] = 5'b00000; w[185][137] = 5'b01111; w[185][138] = 5'b01111; w[185][139] = 5'b01111; w[185][140] = 5'b01111; w[185][141] = 5'b01111; w[185][142] = 5'b01111; w[185][143] = 5'b00000; w[185][144] = 5'b00000; w[185][145] = 5'b01111; w[185][146] = 5'b00000; w[185][147] = 5'b10000; w[185][148] = 5'b01111; w[185][149] = 5'b00000; w[185][150] = 5'b00000; w[185][151] = 5'b01111; w[185][152] = 5'b01111; w[185][153] = 5'b01111; w[185][154] = 5'b01111; w[185][155] = 5'b01111; w[185][156] = 5'b01111; w[185][157] = 5'b00000; w[185][158] = 5'b00000; w[185][159] = 5'b00000; w[185][160] = 5'b10000; w[185][161] = 5'b10000; w[185][162] = 5'b10000; w[185][163] = 5'b00000; w[185][164] = 5'b00000; w[185][165] = 5'b01111; w[185][166] = 5'b01111; w[185][167] = 5'b01111; w[185][168] = 5'b01111; w[185][169] = 5'b01111; w[185][170] = 5'b01111; w[185][171] = 5'b01111; w[185][172] = 5'b00000; w[185][173] = 5'b00000; w[185][174] = 5'b10000; w[185][175] = 5'b10000; w[185][176] = 5'b10000; w[185][177] = 5'b00000; w[185][178] = 5'b01111; w[185][179] = 5'b01111; w[185][180] = 5'b01111; w[185][181] = 5'b01111; w[185][182] = 5'b01111; w[185][183] = 5'b01111; w[185][184] = 5'b01111; w[185][185] = 5'b00000; w[185][186] = 5'b01111; w[185][187] = 5'b01111; w[185][188] = 5'b01111; w[185][189] = 5'b01111; w[185][190] = 5'b01111; w[185][191] = 5'b01111; w[185][192] = 5'b01111; w[185][193] = 5'b01111; w[185][194] = 5'b01111; w[185][195] = 5'b01111; w[185][196] = 5'b01111; w[185][197] = 5'b01111; w[185][198] = 5'b01111; w[185][199] = 5'b01111; w[185][200] = 5'b01111; w[185][201] = 5'b01111; w[185][202] = 5'b01111; w[185][203] = 5'b01111; w[185][204] = 5'b01111; w[185][205] = 5'b01111; w[185][206] = 5'b01111; w[185][207] = 5'b01111; w[185][208] = 5'b01111; w[185][209] = 5'b01111; 
w[186][0] = 5'b01111; w[186][1] = 5'b01111; w[186][2] = 5'b01111; w[186][3] = 5'b01111; w[186][4] = 5'b01111; w[186][5] = 5'b01111; w[186][6] = 5'b01111; w[186][7] = 5'b01111; w[186][8] = 5'b01111; w[186][9] = 5'b01111; w[186][10] = 5'b01111; w[186][11] = 5'b01111; w[186][12] = 5'b01111; w[186][13] = 5'b01111; w[186][14] = 5'b01111; w[186][15] = 5'b01111; w[186][16] = 5'b01111; w[186][17] = 5'b01111; w[186][18] = 5'b01111; w[186][19] = 5'b01111; w[186][20] = 5'b01111; w[186][21] = 5'b01111; w[186][22] = 5'b01111; w[186][23] = 5'b01111; w[186][24] = 5'b01111; w[186][25] = 5'b01111; w[186][26] = 5'b01111; w[186][27] = 5'b01111; w[186][28] = 5'b01111; w[186][29] = 5'b01111; w[186][30] = 5'b01111; w[186][31] = 5'b00000; w[186][32] = 5'b10000; w[186][33] = 5'b10000; w[186][34] = 5'b10000; w[186][35] = 5'b10000; w[186][36] = 5'b10000; w[186][37] = 5'b10000; w[186][38] = 5'b00000; w[186][39] = 5'b01111; w[186][40] = 5'b01111; w[186][41] = 5'b01111; w[186][42] = 5'b01111; w[186][43] = 5'b01111; w[186][44] = 5'b01111; w[186][45] = 5'b10000; w[186][46] = 5'b10000; w[186][47] = 5'b10000; w[186][48] = 5'b10000; w[186][49] = 5'b10000; w[186][50] = 5'b10000; w[186][51] = 5'b10000; w[186][52] = 5'b10000; w[186][53] = 5'b01111; w[186][54] = 5'b01111; w[186][55] = 5'b01111; w[186][56] = 5'b01111; w[186][57] = 5'b01111; w[186][58] = 5'b01111; w[186][59] = 5'b00000; w[186][60] = 5'b00000; w[186][61] = 5'b01111; w[186][62] = 5'b10000; w[186][63] = 5'b00000; w[186][64] = 5'b01111; w[186][65] = 5'b00000; w[186][66] = 5'b00000; w[186][67] = 5'b01111; w[186][68] = 5'b01111; w[186][69] = 5'b01111; w[186][70] = 5'b01111; w[186][71] = 5'b01111; w[186][72] = 5'b01111; w[186][73] = 5'b00000; w[186][74] = 5'b01111; w[186][75] = 5'b01111; w[186][76] = 5'b10000; w[186][77] = 5'b00000; w[186][78] = 5'b01111; w[186][79] = 5'b01111; w[186][80] = 5'b00000; w[186][81] = 5'b01111; w[186][82] = 5'b01111; w[186][83] = 5'b01111; w[186][84] = 5'b01111; w[186][85] = 5'b01111; w[186][86] = 5'b01111; w[186][87] = 5'b00000; w[186][88] = 5'b01111; w[186][89] = 5'b01111; w[186][90] = 5'b10000; w[186][91] = 5'b10000; w[186][92] = 5'b01111; w[186][93] = 5'b01111; w[186][94] = 5'b01111; w[186][95] = 5'b01111; w[186][96] = 5'b01111; w[186][97] = 5'b01111; w[186][98] = 5'b01111; w[186][99] = 5'b01111; w[186][100] = 5'b01111; w[186][101] = 5'b00000; w[186][102] = 5'b01111; w[186][103] = 5'b01111; w[186][104] = 5'b10000; w[186][105] = 5'b10000; w[186][106] = 5'b01111; w[186][107] = 5'b00000; w[186][108] = 5'b00000; w[186][109] = 5'b01111; w[186][110] = 5'b01111; w[186][111] = 5'b01111; w[186][112] = 5'b01111; w[186][113] = 5'b01111; w[186][114] = 5'b01111; w[186][115] = 5'b00000; w[186][116] = 5'b01111; w[186][117] = 5'b01111; w[186][118] = 5'b10000; w[186][119] = 5'b10000; w[186][120] = 5'b00000; w[186][121] = 5'b00000; w[186][122] = 5'b00000; w[186][123] = 5'b01111; w[186][124] = 5'b01111; w[186][125] = 5'b01111; w[186][126] = 5'b01111; w[186][127] = 5'b01111; w[186][128] = 5'b01111; w[186][129] = 5'b00000; w[186][130] = 5'b01111; w[186][131] = 5'b01111; w[186][132] = 5'b00000; w[186][133] = 5'b10000; w[186][134] = 5'b01111; w[186][135] = 5'b01111; w[186][136] = 5'b00000; w[186][137] = 5'b01111; w[186][138] = 5'b01111; w[186][139] = 5'b01111; w[186][140] = 5'b01111; w[186][141] = 5'b01111; w[186][142] = 5'b01111; w[186][143] = 5'b00000; w[186][144] = 5'b00000; w[186][145] = 5'b01111; w[186][146] = 5'b00000; w[186][147] = 5'b10000; w[186][148] = 5'b01111; w[186][149] = 5'b00000; w[186][150] = 5'b00000; w[186][151] = 5'b01111; w[186][152] = 5'b01111; w[186][153] = 5'b01111; w[186][154] = 5'b01111; w[186][155] = 5'b01111; w[186][156] = 5'b01111; w[186][157] = 5'b00000; w[186][158] = 5'b00000; w[186][159] = 5'b00000; w[186][160] = 5'b10000; w[186][161] = 5'b10000; w[186][162] = 5'b10000; w[186][163] = 5'b00000; w[186][164] = 5'b00000; w[186][165] = 5'b01111; w[186][166] = 5'b01111; w[186][167] = 5'b01111; w[186][168] = 5'b01111; w[186][169] = 5'b01111; w[186][170] = 5'b01111; w[186][171] = 5'b01111; w[186][172] = 5'b00000; w[186][173] = 5'b00000; w[186][174] = 5'b10000; w[186][175] = 5'b10000; w[186][176] = 5'b10000; w[186][177] = 5'b00000; w[186][178] = 5'b01111; w[186][179] = 5'b01111; w[186][180] = 5'b01111; w[186][181] = 5'b01111; w[186][182] = 5'b01111; w[186][183] = 5'b01111; w[186][184] = 5'b01111; w[186][185] = 5'b01111; w[186][186] = 5'b00000; w[186][187] = 5'b01111; w[186][188] = 5'b01111; w[186][189] = 5'b01111; w[186][190] = 5'b01111; w[186][191] = 5'b01111; w[186][192] = 5'b01111; w[186][193] = 5'b01111; w[186][194] = 5'b01111; w[186][195] = 5'b01111; w[186][196] = 5'b01111; w[186][197] = 5'b01111; w[186][198] = 5'b01111; w[186][199] = 5'b01111; w[186][200] = 5'b01111; w[186][201] = 5'b01111; w[186][202] = 5'b01111; w[186][203] = 5'b01111; w[186][204] = 5'b01111; w[186][205] = 5'b01111; w[186][206] = 5'b01111; w[186][207] = 5'b01111; w[186][208] = 5'b01111; w[186][209] = 5'b01111; 
w[187][0] = 5'b01111; w[187][1] = 5'b01111; w[187][2] = 5'b01111; w[187][3] = 5'b01111; w[187][4] = 5'b01111; w[187][5] = 5'b01111; w[187][6] = 5'b01111; w[187][7] = 5'b01111; w[187][8] = 5'b01111; w[187][9] = 5'b01111; w[187][10] = 5'b01111; w[187][11] = 5'b01111; w[187][12] = 5'b01111; w[187][13] = 5'b01111; w[187][14] = 5'b01111; w[187][15] = 5'b01111; w[187][16] = 5'b01111; w[187][17] = 5'b01111; w[187][18] = 5'b01111; w[187][19] = 5'b01111; w[187][20] = 5'b01111; w[187][21] = 5'b01111; w[187][22] = 5'b01111; w[187][23] = 5'b01111; w[187][24] = 5'b01111; w[187][25] = 5'b01111; w[187][26] = 5'b01111; w[187][27] = 5'b01111; w[187][28] = 5'b01111; w[187][29] = 5'b01111; w[187][30] = 5'b01111; w[187][31] = 5'b00000; w[187][32] = 5'b10000; w[187][33] = 5'b10000; w[187][34] = 5'b10000; w[187][35] = 5'b10000; w[187][36] = 5'b10000; w[187][37] = 5'b10000; w[187][38] = 5'b00000; w[187][39] = 5'b01111; w[187][40] = 5'b01111; w[187][41] = 5'b01111; w[187][42] = 5'b01111; w[187][43] = 5'b01111; w[187][44] = 5'b01111; w[187][45] = 5'b10000; w[187][46] = 5'b10000; w[187][47] = 5'b10000; w[187][48] = 5'b10000; w[187][49] = 5'b10000; w[187][50] = 5'b10000; w[187][51] = 5'b10000; w[187][52] = 5'b10000; w[187][53] = 5'b01111; w[187][54] = 5'b01111; w[187][55] = 5'b01111; w[187][56] = 5'b01111; w[187][57] = 5'b01111; w[187][58] = 5'b01111; w[187][59] = 5'b00000; w[187][60] = 5'b00000; w[187][61] = 5'b01111; w[187][62] = 5'b10000; w[187][63] = 5'b00000; w[187][64] = 5'b01111; w[187][65] = 5'b00000; w[187][66] = 5'b00000; w[187][67] = 5'b01111; w[187][68] = 5'b01111; w[187][69] = 5'b01111; w[187][70] = 5'b01111; w[187][71] = 5'b01111; w[187][72] = 5'b01111; w[187][73] = 5'b00000; w[187][74] = 5'b01111; w[187][75] = 5'b01111; w[187][76] = 5'b10000; w[187][77] = 5'b00000; w[187][78] = 5'b01111; w[187][79] = 5'b01111; w[187][80] = 5'b00000; w[187][81] = 5'b01111; w[187][82] = 5'b01111; w[187][83] = 5'b01111; w[187][84] = 5'b01111; w[187][85] = 5'b01111; w[187][86] = 5'b01111; w[187][87] = 5'b00000; w[187][88] = 5'b01111; w[187][89] = 5'b01111; w[187][90] = 5'b10000; w[187][91] = 5'b10000; w[187][92] = 5'b01111; w[187][93] = 5'b01111; w[187][94] = 5'b01111; w[187][95] = 5'b01111; w[187][96] = 5'b01111; w[187][97] = 5'b01111; w[187][98] = 5'b01111; w[187][99] = 5'b01111; w[187][100] = 5'b01111; w[187][101] = 5'b00000; w[187][102] = 5'b01111; w[187][103] = 5'b01111; w[187][104] = 5'b10000; w[187][105] = 5'b10000; w[187][106] = 5'b01111; w[187][107] = 5'b00000; w[187][108] = 5'b00000; w[187][109] = 5'b01111; w[187][110] = 5'b01111; w[187][111] = 5'b01111; w[187][112] = 5'b01111; w[187][113] = 5'b01111; w[187][114] = 5'b01111; w[187][115] = 5'b00000; w[187][116] = 5'b01111; w[187][117] = 5'b01111; w[187][118] = 5'b10000; w[187][119] = 5'b10000; w[187][120] = 5'b00000; w[187][121] = 5'b00000; w[187][122] = 5'b00000; w[187][123] = 5'b01111; w[187][124] = 5'b01111; w[187][125] = 5'b01111; w[187][126] = 5'b01111; w[187][127] = 5'b01111; w[187][128] = 5'b01111; w[187][129] = 5'b00000; w[187][130] = 5'b01111; w[187][131] = 5'b01111; w[187][132] = 5'b00000; w[187][133] = 5'b10000; w[187][134] = 5'b01111; w[187][135] = 5'b01111; w[187][136] = 5'b00000; w[187][137] = 5'b01111; w[187][138] = 5'b01111; w[187][139] = 5'b01111; w[187][140] = 5'b01111; w[187][141] = 5'b01111; w[187][142] = 5'b01111; w[187][143] = 5'b00000; w[187][144] = 5'b00000; w[187][145] = 5'b01111; w[187][146] = 5'b00000; w[187][147] = 5'b10000; w[187][148] = 5'b01111; w[187][149] = 5'b00000; w[187][150] = 5'b00000; w[187][151] = 5'b01111; w[187][152] = 5'b01111; w[187][153] = 5'b01111; w[187][154] = 5'b01111; w[187][155] = 5'b01111; w[187][156] = 5'b01111; w[187][157] = 5'b00000; w[187][158] = 5'b00000; w[187][159] = 5'b00000; w[187][160] = 5'b10000; w[187][161] = 5'b10000; w[187][162] = 5'b10000; w[187][163] = 5'b00000; w[187][164] = 5'b00000; w[187][165] = 5'b01111; w[187][166] = 5'b01111; w[187][167] = 5'b01111; w[187][168] = 5'b01111; w[187][169] = 5'b01111; w[187][170] = 5'b01111; w[187][171] = 5'b01111; w[187][172] = 5'b00000; w[187][173] = 5'b00000; w[187][174] = 5'b10000; w[187][175] = 5'b10000; w[187][176] = 5'b10000; w[187][177] = 5'b00000; w[187][178] = 5'b01111; w[187][179] = 5'b01111; w[187][180] = 5'b01111; w[187][181] = 5'b01111; w[187][182] = 5'b01111; w[187][183] = 5'b01111; w[187][184] = 5'b01111; w[187][185] = 5'b01111; w[187][186] = 5'b01111; w[187][187] = 5'b00000; w[187][188] = 5'b01111; w[187][189] = 5'b01111; w[187][190] = 5'b01111; w[187][191] = 5'b01111; w[187][192] = 5'b01111; w[187][193] = 5'b01111; w[187][194] = 5'b01111; w[187][195] = 5'b01111; w[187][196] = 5'b01111; w[187][197] = 5'b01111; w[187][198] = 5'b01111; w[187][199] = 5'b01111; w[187][200] = 5'b01111; w[187][201] = 5'b01111; w[187][202] = 5'b01111; w[187][203] = 5'b01111; w[187][204] = 5'b01111; w[187][205] = 5'b01111; w[187][206] = 5'b01111; w[187][207] = 5'b01111; w[187][208] = 5'b01111; w[187][209] = 5'b01111; 
w[188][0] = 5'b01111; w[188][1] = 5'b01111; w[188][2] = 5'b01111; w[188][3] = 5'b01111; w[188][4] = 5'b01111; w[188][5] = 5'b01111; w[188][6] = 5'b01111; w[188][7] = 5'b01111; w[188][8] = 5'b01111; w[188][9] = 5'b01111; w[188][10] = 5'b01111; w[188][11] = 5'b01111; w[188][12] = 5'b01111; w[188][13] = 5'b01111; w[188][14] = 5'b01111; w[188][15] = 5'b01111; w[188][16] = 5'b01111; w[188][17] = 5'b01111; w[188][18] = 5'b01111; w[188][19] = 5'b01111; w[188][20] = 5'b01111; w[188][21] = 5'b01111; w[188][22] = 5'b01111; w[188][23] = 5'b01111; w[188][24] = 5'b01111; w[188][25] = 5'b01111; w[188][26] = 5'b01111; w[188][27] = 5'b01111; w[188][28] = 5'b01111; w[188][29] = 5'b01111; w[188][30] = 5'b01111; w[188][31] = 5'b00000; w[188][32] = 5'b10000; w[188][33] = 5'b10000; w[188][34] = 5'b10000; w[188][35] = 5'b10000; w[188][36] = 5'b10000; w[188][37] = 5'b10000; w[188][38] = 5'b00000; w[188][39] = 5'b01111; w[188][40] = 5'b01111; w[188][41] = 5'b01111; w[188][42] = 5'b01111; w[188][43] = 5'b01111; w[188][44] = 5'b01111; w[188][45] = 5'b10000; w[188][46] = 5'b10000; w[188][47] = 5'b10000; w[188][48] = 5'b10000; w[188][49] = 5'b10000; w[188][50] = 5'b10000; w[188][51] = 5'b10000; w[188][52] = 5'b10000; w[188][53] = 5'b01111; w[188][54] = 5'b01111; w[188][55] = 5'b01111; w[188][56] = 5'b01111; w[188][57] = 5'b01111; w[188][58] = 5'b01111; w[188][59] = 5'b00000; w[188][60] = 5'b00000; w[188][61] = 5'b01111; w[188][62] = 5'b10000; w[188][63] = 5'b00000; w[188][64] = 5'b01111; w[188][65] = 5'b00000; w[188][66] = 5'b00000; w[188][67] = 5'b01111; w[188][68] = 5'b01111; w[188][69] = 5'b01111; w[188][70] = 5'b01111; w[188][71] = 5'b01111; w[188][72] = 5'b01111; w[188][73] = 5'b00000; w[188][74] = 5'b01111; w[188][75] = 5'b01111; w[188][76] = 5'b10000; w[188][77] = 5'b00000; w[188][78] = 5'b01111; w[188][79] = 5'b01111; w[188][80] = 5'b00000; w[188][81] = 5'b01111; w[188][82] = 5'b01111; w[188][83] = 5'b01111; w[188][84] = 5'b01111; w[188][85] = 5'b01111; w[188][86] = 5'b01111; w[188][87] = 5'b00000; w[188][88] = 5'b01111; w[188][89] = 5'b01111; w[188][90] = 5'b10000; w[188][91] = 5'b10000; w[188][92] = 5'b01111; w[188][93] = 5'b01111; w[188][94] = 5'b01111; w[188][95] = 5'b01111; w[188][96] = 5'b01111; w[188][97] = 5'b01111; w[188][98] = 5'b01111; w[188][99] = 5'b01111; w[188][100] = 5'b01111; w[188][101] = 5'b00000; w[188][102] = 5'b01111; w[188][103] = 5'b01111; w[188][104] = 5'b10000; w[188][105] = 5'b10000; w[188][106] = 5'b01111; w[188][107] = 5'b00000; w[188][108] = 5'b00000; w[188][109] = 5'b01111; w[188][110] = 5'b01111; w[188][111] = 5'b01111; w[188][112] = 5'b01111; w[188][113] = 5'b01111; w[188][114] = 5'b01111; w[188][115] = 5'b00000; w[188][116] = 5'b01111; w[188][117] = 5'b01111; w[188][118] = 5'b10000; w[188][119] = 5'b10000; w[188][120] = 5'b00000; w[188][121] = 5'b00000; w[188][122] = 5'b00000; w[188][123] = 5'b01111; w[188][124] = 5'b01111; w[188][125] = 5'b01111; w[188][126] = 5'b01111; w[188][127] = 5'b01111; w[188][128] = 5'b01111; w[188][129] = 5'b00000; w[188][130] = 5'b01111; w[188][131] = 5'b01111; w[188][132] = 5'b00000; w[188][133] = 5'b10000; w[188][134] = 5'b01111; w[188][135] = 5'b01111; w[188][136] = 5'b00000; w[188][137] = 5'b01111; w[188][138] = 5'b01111; w[188][139] = 5'b01111; w[188][140] = 5'b01111; w[188][141] = 5'b01111; w[188][142] = 5'b01111; w[188][143] = 5'b00000; w[188][144] = 5'b00000; w[188][145] = 5'b01111; w[188][146] = 5'b00000; w[188][147] = 5'b10000; w[188][148] = 5'b01111; w[188][149] = 5'b00000; w[188][150] = 5'b00000; w[188][151] = 5'b01111; w[188][152] = 5'b01111; w[188][153] = 5'b01111; w[188][154] = 5'b01111; w[188][155] = 5'b01111; w[188][156] = 5'b01111; w[188][157] = 5'b00000; w[188][158] = 5'b00000; w[188][159] = 5'b00000; w[188][160] = 5'b10000; w[188][161] = 5'b10000; w[188][162] = 5'b10000; w[188][163] = 5'b00000; w[188][164] = 5'b00000; w[188][165] = 5'b01111; w[188][166] = 5'b01111; w[188][167] = 5'b01111; w[188][168] = 5'b01111; w[188][169] = 5'b01111; w[188][170] = 5'b01111; w[188][171] = 5'b01111; w[188][172] = 5'b00000; w[188][173] = 5'b00000; w[188][174] = 5'b10000; w[188][175] = 5'b10000; w[188][176] = 5'b10000; w[188][177] = 5'b00000; w[188][178] = 5'b01111; w[188][179] = 5'b01111; w[188][180] = 5'b01111; w[188][181] = 5'b01111; w[188][182] = 5'b01111; w[188][183] = 5'b01111; w[188][184] = 5'b01111; w[188][185] = 5'b01111; w[188][186] = 5'b01111; w[188][187] = 5'b01111; w[188][188] = 5'b00000; w[188][189] = 5'b01111; w[188][190] = 5'b01111; w[188][191] = 5'b01111; w[188][192] = 5'b01111; w[188][193] = 5'b01111; w[188][194] = 5'b01111; w[188][195] = 5'b01111; w[188][196] = 5'b01111; w[188][197] = 5'b01111; w[188][198] = 5'b01111; w[188][199] = 5'b01111; w[188][200] = 5'b01111; w[188][201] = 5'b01111; w[188][202] = 5'b01111; w[188][203] = 5'b01111; w[188][204] = 5'b01111; w[188][205] = 5'b01111; w[188][206] = 5'b01111; w[188][207] = 5'b01111; w[188][208] = 5'b01111; w[188][209] = 5'b01111; 
w[189][0] = 5'b01111; w[189][1] = 5'b01111; w[189][2] = 5'b01111; w[189][3] = 5'b01111; w[189][4] = 5'b01111; w[189][5] = 5'b01111; w[189][6] = 5'b01111; w[189][7] = 5'b01111; w[189][8] = 5'b01111; w[189][9] = 5'b01111; w[189][10] = 5'b01111; w[189][11] = 5'b01111; w[189][12] = 5'b01111; w[189][13] = 5'b01111; w[189][14] = 5'b01111; w[189][15] = 5'b01111; w[189][16] = 5'b01111; w[189][17] = 5'b01111; w[189][18] = 5'b01111; w[189][19] = 5'b01111; w[189][20] = 5'b01111; w[189][21] = 5'b01111; w[189][22] = 5'b01111; w[189][23] = 5'b01111; w[189][24] = 5'b01111; w[189][25] = 5'b01111; w[189][26] = 5'b01111; w[189][27] = 5'b01111; w[189][28] = 5'b01111; w[189][29] = 5'b01111; w[189][30] = 5'b01111; w[189][31] = 5'b00000; w[189][32] = 5'b10000; w[189][33] = 5'b10000; w[189][34] = 5'b10000; w[189][35] = 5'b10000; w[189][36] = 5'b10000; w[189][37] = 5'b10000; w[189][38] = 5'b00000; w[189][39] = 5'b01111; w[189][40] = 5'b01111; w[189][41] = 5'b01111; w[189][42] = 5'b01111; w[189][43] = 5'b01111; w[189][44] = 5'b01111; w[189][45] = 5'b10000; w[189][46] = 5'b10000; w[189][47] = 5'b10000; w[189][48] = 5'b10000; w[189][49] = 5'b10000; w[189][50] = 5'b10000; w[189][51] = 5'b10000; w[189][52] = 5'b10000; w[189][53] = 5'b01111; w[189][54] = 5'b01111; w[189][55] = 5'b01111; w[189][56] = 5'b01111; w[189][57] = 5'b01111; w[189][58] = 5'b01111; w[189][59] = 5'b00000; w[189][60] = 5'b00000; w[189][61] = 5'b01111; w[189][62] = 5'b10000; w[189][63] = 5'b00000; w[189][64] = 5'b01111; w[189][65] = 5'b00000; w[189][66] = 5'b00000; w[189][67] = 5'b01111; w[189][68] = 5'b01111; w[189][69] = 5'b01111; w[189][70] = 5'b01111; w[189][71] = 5'b01111; w[189][72] = 5'b01111; w[189][73] = 5'b00000; w[189][74] = 5'b01111; w[189][75] = 5'b01111; w[189][76] = 5'b10000; w[189][77] = 5'b00000; w[189][78] = 5'b01111; w[189][79] = 5'b01111; w[189][80] = 5'b00000; w[189][81] = 5'b01111; w[189][82] = 5'b01111; w[189][83] = 5'b01111; w[189][84] = 5'b01111; w[189][85] = 5'b01111; w[189][86] = 5'b01111; w[189][87] = 5'b00000; w[189][88] = 5'b01111; w[189][89] = 5'b01111; w[189][90] = 5'b10000; w[189][91] = 5'b10000; w[189][92] = 5'b01111; w[189][93] = 5'b01111; w[189][94] = 5'b01111; w[189][95] = 5'b01111; w[189][96] = 5'b01111; w[189][97] = 5'b01111; w[189][98] = 5'b01111; w[189][99] = 5'b01111; w[189][100] = 5'b01111; w[189][101] = 5'b00000; w[189][102] = 5'b01111; w[189][103] = 5'b01111; w[189][104] = 5'b10000; w[189][105] = 5'b10000; w[189][106] = 5'b01111; w[189][107] = 5'b00000; w[189][108] = 5'b00000; w[189][109] = 5'b01111; w[189][110] = 5'b01111; w[189][111] = 5'b01111; w[189][112] = 5'b01111; w[189][113] = 5'b01111; w[189][114] = 5'b01111; w[189][115] = 5'b00000; w[189][116] = 5'b01111; w[189][117] = 5'b01111; w[189][118] = 5'b10000; w[189][119] = 5'b10000; w[189][120] = 5'b00000; w[189][121] = 5'b00000; w[189][122] = 5'b00000; w[189][123] = 5'b01111; w[189][124] = 5'b01111; w[189][125] = 5'b01111; w[189][126] = 5'b01111; w[189][127] = 5'b01111; w[189][128] = 5'b01111; w[189][129] = 5'b00000; w[189][130] = 5'b01111; w[189][131] = 5'b01111; w[189][132] = 5'b00000; w[189][133] = 5'b10000; w[189][134] = 5'b01111; w[189][135] = 5'b01111; w[189][136] = 5'b00000; w[189][137] = 5'b01111; w[189][138] = 5'b01111; w[189][139] = 5'b01111; w[189][140] = 5'b01111; w[189][141] = 5'b01111; w[189][142] = 5'b01111; w[189][143] = 5'b00000; w[189][144] = 5'b00000; w[189][145] = 5'b01111; w[189][146] = 5'b00000; w[189][147] = 5'b10000; w[189][148] = 5'b01111; w[189][149] = 5'b00000; w[189][150] = 5'b00000; w[189][151] = 5'b01111; w[189][152] = 5'b01111; w[189][153] = 5'b01111; w[189][154] = 5'b01111; w[189][155] = 5'b01111; w[189][156] = 5'b01111; w[189][157] = 5'b00000; w[189][158] = 5'b00000; w[189][159] = 5'b00000; w[189][160] = 5'b10000; w[189][161] = 5'b10000; w[189][162] = 5'b10000; w[189][163] = 5'b00000; w[189][164] = 5'b00000; w[189][165] = 5'b01111; w[189][166] = 5'b01111; w[189][167] = 5'b01111; w[189][168] = 5'b01111; w[189][169] = 5'b01111; w[189][170] = 5'b01111; w[189][171] = 5'b01111; w[189][172] = 5'b00000; w[189][173] = 5'b00000; w[189][174] = 5'b10000; w[189][175] = 5'b10000; w[189][176] = 5'b10000; w[189][177] = 5'b00000; w[189][178] = 5'b01111; w[189][179] = 5'b01111; w[189][180] = 5'b01111; w[189][181] = 5'b01111; w[189][182] = 5'b01111; w[189][183] = 5'b01111; w[189][184] = 5'b01111; w[189][185] = 5'b01111; w[189][186] = 5'b01111; w[189][187] = 5'b01111; w[189][188] = 5'b01111; w[189][189] = 5'b00000; w[189][190] = 5'b01111; w[189][191] = 5'b01111; w[189][192] = 5'b01111; w[189][193] = 5'b01111; w[189][194] = 5'b01111; w[189][195] = 5'b01111; w[189][196] = 5'b01111; w[189][197] = 5'b01111; w[189][198] = 5'b01111; w[189][199] = 5'b01111; w[189][200] = 5'b01111; w[189][201] = 5'b01111; w[189][202] = 5'b01111; w[189][203] = 5'b01111; w[189][204] = 5'b01111; w[189][205] = 5'b01111; w[189][206] = 5'b01111; w[189][207] = 5'b01111; w[189][208] = 5'b01111; w[189][209] = 5'b01111; 
w[190][0] = 5'b01111; w[190][1] = 5'b01111; w[190][2] = 5'b01111; w[190][3] = 5'b01111; w[190][4] = 5'b01111; w[190][5] = 5'b01111; w[190][6] = 5'b01111; w[190][7] = 5'b01111; w[190][8] = 5'b01111; w[190][9] = 5'b01111; w[190][10] = 5'b01111; w[190][11] = 5'b01111; w[190][12] = 5'b01111; w[190][13] = 5'b01111; w[190][14] = 5'b01111; w[190][15] = 5'b01111; w[190][16] = 5'b01111; w[190][17] = 5'b01111; w[190][18] = 5'b01111; w[190][19] = 5'b01111; w[190][20] = 5'b01111; w[190][21] = 5'b01111; w[190][22] = 5'b01111; w[190][23] = 5'b01111; w[190][24] = 5'b01111; w[190][25] = 5'b01111; w[190][26] = 5'b01111; w[190][27] = 5'b01111; w[190][28] = 5'b01111; w[190][29] = 5'b01111; w[190][30] = 5'b01111; w[190][31] = 5'b00000; w[190][32] = 5'b10000; w[190][33] = 5'b10000; w[190][34] = 5'b10000; w[190][35] = 5'b10000; w[190][36] = 5'b10000; w[190][37] = 5'b10000; w[190][38] = 5'b00000; w[190][39] = 5'b01111; w[190][40] = 5'b01111; w[190][41] = 5'b01111; w[190][42] = 5'b01111; w[190][43] = 5'b01111; w[190][44] = 5'b01111; w[190][45] = 5'b10000; w[190][46] = 5'b10000; w[190][47] = 5'b10000; w[190][48] = 5'b10000; w[190][49] = 5'b10000; w[190][50] = 5'b10000; w[190][51] = 5'b10000; w[190][52] = 5'b10000; w[190][53] = 5'b01111; w[190][54] = 5'b01111; w[190][55] = 5'b01111; w[190][56] = 5'b01111; w[190][57] = 5'b01111; w[190][58] = 5'b01111; w[190][59] = 5'b00000; w[190][60] = 5'b00000; w[190][61] = 5'b01111; w[190][62] = 5'b10000; w[190][63] = 5'b00000; w[190][64] = 5'b01111; w[190][65] = 5'b00000; w[190][66] = 5'b00000; w[190][67] = 5'b01111; w[190][68] = 5'b01111; w[190][69] = 5'b01111; w[190][70] = 5'b01111; w[190][71] = 5'b01111; w[190][72] = 5'b01111; w[190][73] = 5'b00000; w[190][74] = 5'b01111; w[190][75] = 5'b01111; w[190][76] = 5'b10000; w[190][77] = 5'b00000; w[190][78] = 5'b01111; w[190][79] = 5'b01111; w[190][80] = 5'b00000; w[190][81] = 5'b01111; w[190][82] = 5'b01111; w[190][83] = 5'b01111; w[190][84] = 5'b01111; w[190][85] = 5'b01111; w[190][86] = 5'b01111; w[190][87] = 5'b00000; w[190][88] = 5'b01111; w[190][89] = 5'b01111; w[190][90] = 5'b10000; w[190][91] = 5'b10000; w[190][92] = 5'b01111; w[190][93] = 5'b01111; w[190][94] = 5'b01111; w[190][95] = 5'b01111; w[190][96] = 5'b01111; w[190][97] = 5'b01111; w[190][98] = 5'b01111; w[190][99] = 5'b01111; w[190][100] = 5'b01111; w[190][101] = 5'b00000; w[190][102] = 5'b01111; w[190][103] = 5'b01111; w[190][104] = 5'b10000; w[190][105] = 5'b10000; w[190][106] = 5'b01111; w[190][107] = 5'b00000; w[190][108] = 5'b00000; w[190][109] = 5'b01111; w[190][110] = 5'b01111; w[190][111] = 5'b01111; w[190][112] = 5'b01111; w[190][113] = 5'b01111; w[190][114] = 5'b01111; w[190][115] = 5'b00000; w[190][116] = 5'b01111; w[190][117] = 5'b01111; w[190][118] = 5'b10000; w[190][119] = 5'b10000; w[190][120] = 5'b00000; w[190][121] = 5'b00000; w[190][122] = 5'b00000; w[190][123] = 5'b01111; w[190][124] = 5'b01111; w[190][125] = 5'b01111; w[190][126] = 5'b01111; w[190][127] = 5'b01111; w[190][128] = 5'b01111; w[190][129] = 5'b00000; w[190][130] = 5'b01111; w[190][131] = 5'b01111; w[190][132] = 5'b00000; w[190][133] = 5'b10000; w[190][134] = 5'b01111; w[190][135] = 5'b01111; w[190][136] = 5'b00000; w[190][137] = 5'b01111; w[190][138] = 5'b01111; w[190][139] = 5'b01111; w[190][140] = 5'b01111; w[190][141] = 5'b01111; w[190][142] = 5'b01111; w[190][143] = 5'b00000; w[190][144] = 5'b00000; w[190][145] = 5'b01111; w[190][146] = 5'b00000; w[190][147] = 5'b10000; w[190][148] = 5'b01111; w[190][149] = 5'b00000; w[190][150] = 5'b00000; w[190][151] = 5'b01111; w[190][152] = 5'b01111; w[190][153] = 5'b01111; w[190][154] = 5'b01111; w[190][155] = 5'b01111; w[190][156] = 5'b01111; w[190][157] = 5'b00000; w[190][158] = 5'b00000; w[190][159] = 5'b00000; w[190][160] = 5'b10000; w[190][161] = 5'b10000; w[190][162] = 5'b10000; w[190][163] = 5'b00000; w[190][164] = 5'b00000; w[190][165] = 5'b01111; w[190][166] = 5'b01111; w[190][167] = 5'b01111; w[190][168] = 5'b01111; w[190][169] = 5'b01111; w[190][170] = 5'b01111; w[190][171] = 5'b01111; w[190][172] = 5'b00000; w[190][173] = 5'b00000; w[190][174] = 5'b10000; w[190][175] = 5'b10000; w[190][176] = 5'b10000; w[190][177] = 5'b00000; w[190][178] = 5'b01111; w[190][179] = 5'b01111; w[190][180] = 5'b01111; w[190][181] = 5'b01111; w[190][182] = 5'b01111; w[190][183] = 5'b01111; w[190][184] = 5'b01111; w[190][185] = 5'b01111; w[190][186] = 5'b01111; w[190][187] = 5'b01111; w[190][188] = 5'b01111; w[190][189] = 5'b01111; w[190][190] = 5'b00000; w[190][191] = 5'b01111; w[190][192] = 5'b01111; w[190][193] = 5'b01111; w[190][194] = 5'b01111; w[190][195] = 5'b01111; w[190][196] = 5'b01111; w[190][197] = 5'b01111; w[190][198] = 5'b01111; w[190][199] = 5'b01111; w[190][200] = 5'b01111; w[190][201] = 5'b01111; w[190][202] = 5'b01111; w[190][203] = 5'b01111; w[190][204] = 5'b01111; w[190][205] = 5'b01111; w[190][206] = 5'b01111; w[190][207] = 5'b01111; w[190][208] = 5'b01111; w[190][209] = 5'b01111; 
w[191][0] = 5'b01111; w[191][1] = 5'b01111; w[191][2] = 5'b01111; w[191][3] = 5'b01111; w[191][4] = 5'b01111; w[191][5] = 5'b01111; w[191][6] = 5'b01111; w[191][7] = 5'b01111; w[191][8] = 5'b01111; w[191][9] = 5'b01111; w[191][10] = 5'b01111; w[191][11] = 5'b01111; w[191][12] = 5'b01111; w[191][13] = 5'b01111; w[191][14] = 5'b01111; w[191][15] = 5'b01111; w[191][16] = 5'b01111; w[191][17] = 5'b01111; w[191][18] = 5'b01111; w[191][19] = 5'b01111; w[191][20] = 5'b01111; w[191][21] = 5'b01111; w[191][22] = 5'b01111; w[191][23] = 5'b01111; w[191][24] = 5'b01111; w[191][25] = 5'b01111; w[191][26] = 5'b01111; w[191][27] = 5'b01111; w[191][28] = 5'b01111; w[191][29] = 5'b01111; w[191][30] = 5'b01111; w[191][31] = 5'b00000; w[191][32] = 5'b10000; w[191][33] = 5'b10000; w[191][34] = 5'b10000; w[191][35] = 5'b10000; w[191][36] = 5'b10000; w[191][37] = 5'b10000; w[191][38] = 5'b00000; w[191][39] = 5'b01111; w[191][40] = 5'b01111; w[191][41] = 5'b01111; w[191][42] = 5'b01111; w[191][43] = 5'b01111; w[191][44] = 5'b01111; w[191][45] = 5'b10000; w[191][46] = 5'b10000; w[191][47] = 5'b10000; w[191][48] = 5'b10000; w[191][49] = 5'b10000; w[191][50] = 5'b10000; w[191][51] = 5'b10000; w[191][52] = 5'b10000; w[191][53] = 5'b01111; w[191][54] = 5'b01111; w[191][55] = 5'b01111; w[191][56] = 5'b01111; w[191][57] = 5'b01111; w[191][58] = 5'b01111; w[191][59] = 5'b00000; w[191][60] = 5'b00000; w[191][61] = 5'b01111; w[191][62] = 5'b10000; w[191][63] = 5'b00000; w[191][64] = 5'b01111; w[191][65] = 5'b00000; w[191][66] = 5'b00000; w[191][67] = 5'b01111; w[191][68] = 5'b01111; w[191][69] = 5'b01111; w[191][70] = 5'b01111; w[191][71] = 5'b01111; w[191][72] = 5'b01111; w[191][73] = 5'b00000; w[191][74] = 5'b01111; w[191][75] = 5'b01111; w[191][76] = 5'b10000; w[191][77] = 5'b00000; w[191][78] = 5'b01111; w[191][79] = 5'b01111; w[191][80] = 5'b00000; w[191][81] = 5'b01111; w[191][82] = 5'b01111; w[191][83] = 5'b01111; w[191][84] = 5'b01111; w[191][85] = 5'b01111; w[191][86] = 5'b01111; w[191][87] = 5'b00000; w[191][88] = 5'b01111; w[191][89] = 5'b01111; w[191][90] = 5'b10000; w[191][91] = 5'b10000; w[191][92] = 5'b01111; w[191][93] = 5'b01111; w[191][94] = 5'b01111; w[191][95] = 5'b01111; w[191][96] = 5'b01111; w[191][97] = 5'b01111; w[191][98] = 5'b01111; w[191][99] = 5'b01111; w[191][100] = 5'b01111; w[191][101] = 5'b00000; w[191][102] = 5'b01111; w[191][103] = 5'b01111; w[191][104] = 5'b10000; w[191][105] = 5'b10000; w[191][106] = 5'b01111; w[191][107] = 5'b00000; w[191][108] = 5'b00000; w[191][109] = 5'b01111; w[191][110] = 5'b01111; w[191][111] = 5'b01111; w[191][112] = 5'b01111; w[191][113] = 5'b01111; w[191][114] = 5'b01111; w[191][115] = 5'b00000; w[191][116] = 5'b01111; w[191][117] = 5'b01111; w[191][118] = 5'b10000; w[191][119] = 5'b10000; w[191][120] = 5'b00000; w[191][121] = 5'b00000; w[191][122] = 5'b00000; w[191][123] = 5'b01111; w[191][124] = 5'b01111; w[191][125] = 5'b01111; w[191][126] = 5'b01111; w[191][127] = 5'b01111; w[191][128] = 5'b01111; w[191][129] = 5'b00000; w[191][130] = 5'b01111; w[191][131] = 5'b01111; w[191][132] = 5'b00000; w[191][133] = 5'b10000; w[191][134] = 5'b01111; w[191][135] = 5'b01111; w[191][136] = 5'b00000; w[191][137] = 5'b01111; w[191][138] = 5'b01111; w[191][139] = 5'b01111; w[191][140] = 5'b01111; w[191][141] = 5'b01111; w[191][142] = 5'b01111; w[191][143] = 5'b00000; w[191][144] = 5'b00000; w[191][145] = 5'b01111; w[191][146] = 5'b00000; w[191][147] = 5'b10000; w[191][148] = 5'b01111; w[191][149] = 5'b00000; w[191][150] = 5'b00000; w[191][151] = 5'b01111; w[191][152] = 5'b01111; w[191][153] = 5'b01111; w[191][154] = 5'b01111; w[191][155] = 5'b01111; w[191][156] = 5'b01111; w[191][157] = 5'b00000; w[191][158] = 5'b00000; w[191][159] = 5'b00000; w[191][160] = 5'b10000; w[191][161] = 5'b10000; w[191][162] = 5'b10000; w[191][163] = 5'b00000; w[191][164] = 5'b00000; w[191][165] = 5'b01111; w[191][166] = 5'b01111; w[191][167] = 5'b01111; w[191][168] = 5'b01111; w[191][169] = 5'b01111; w[191][170] = 5'b01111; w[191][171] = 5'b01111; w[191][172] = 5'b00000; w[191][173] = 5'b00000; w[191][174] = 5'b10000; w[191][175] = 5'b10000; w[191][176] = 5'b10000; w[191][177] = 5'b00000; w[191][178] = 5'b01111; w[191][179] = 5'b01111; w[191][180] = 5'b01111; w[191][181] = 5'b01111; w[191][182] = 5'b01111; w[191][183] = 5'b01111; w[191][184] = 5'b01111; w[191][185] = 5'b01111; w[191][186] = 5'b01111; w[191][187] = 5'b01111; w[191][188] = 5'b01111; w[191][189] = 5'b01111; w[191][190] = 5'b01111; w[191][191] = 5'b00000; w[191][192] = 5'b01111; w[191][193] = 5'b01111; w[191][194] = 5'b01111; w[191][195] = 5'b01111; w[191][196] = 5'b01111; w[191][197] = 5'b01111; w[191][198] = 5'b01111; w[191][199] = 5'b01111; w[191][200] = 5'b01111; w[191][201] = 5'b01111; w[191][202] = 5'b01111; w[191][203] = 5'b01111; w[191][204] = 5'b01111; w[191][205] = 5'b01111; w[191][206] = 5'b01111; w[191][207] = 5'b01111; w[191][208] = 5'b01111; w[191][209] = 5'b01111; 
w[192][0] = 5'b01111; w[192][1] = 5'b01111; w[192][2] = 5'b01111; w[192][3] = 5'b01111; w[192][4] = 5'b01111; w[192][5] = 5'b01111; w[192][6] = 5'b01111; w[192][7] = 5'b01111; w[192][8] = 5'b01111; w[192][9] = 5'b01111; w[192][10] = 5'b01111; w[192][11] = 5'b01111; w[192][12] = 5'b01111; w[192][13] = 5'b01111; w[192][14] = 5'b01111; w[192][15] = 5'b01111; w[192][16] = 5'b01111; w[192][17] = 5'b01111; w[192][18] = 5'b01111; w[192][19] = 5'b01111; w[192][20] = 5'b01111; w[192][21] = 5'b01111; w[192][22] = 5'b01111; w[192][23] = 5'b01111; w[192][24] = 5'b01111; w[192][25] = 5'b01111; w[192][26] = 5'b01111; w[192][27] = 5'b01111; w[192][28] = 5'b01111; w[192][29] = 5'b01111; w[192][30] = 5'b01111; w[192][31] = 5'b00000; w[192][32] = 5'b10000; w[192][33] = 5'b10000; w[192][34] = 5'b10000; w[192][35] = 5'b10000; w[192][36] = 5'b10000; w[192][37] = 5'b10000; w[192][38] = 5'b00000; w[192][39] = 5'b01111; w[192][40] = 5'b01111; w[192][41] = 5'b01111; w[192][42] = 5'b01111; w[192][43] = 5'b01111; w[192][44] = 5'b01111; w[192][45] = 5'b10000; w[192][46] = 5'b10000; w[192][47] = 5'b10000; w[192][48] = 5'b10000; w[192][49] = 5'b10000; w[192][50] = 5'b10000; w[192][51] = 5'b10000; w[192][52] = 5'b10000; w[192][53] = 5'b01111; w[192][54] = 5'b01111; w[192][55] = 5'b01111; w[192][56] = 5'b01111; w[192][57] = 5'b01111; w[192][58] = 5'b01111; w[192][59] = 5'b00000; w[192][60] = 5'b00000; w[192][61] = 5'b01111; w[192][62] = 5'b10000; w[192][63] = 5'b00000; w[192][64] = 5'b01111; w[192][65] = 5'b00000; w[192][66] = 5'b00000; w[192][67] = 5'b01111; w[192][68] = 5'b01111; w[192][69] = 5'b01111; w[192][70] = 5'b01111; w[192][71] = 5'b01111; w[192][72] = 5'b01111; w[192][73] = 5'b00000; w[192][74] = 5'b01111; w[192][75] = 5'b01111; w[192][76] = 5'b10000; w[192][77] = 5'b00000; w[192][78] = 5'b01111; w[192][79] = 5'b01111; w[192][80] = 5'b00000; w[192][81] = 5'b01111; w[192][82] = 5'b01111; w[192][83] = 5'b01111; w[192][84] = 5'b01111; w[192][85] = 5'b01111; w[192][86] = 5'b01111; w[192][87] = 5'b00000; w[192][88] = 5'b01111; w[192][89] = 5'b01111; w[192][90] = 5'b10000; w[192][91] = 5'b10000; w[192][92] = 5'b01111; w[192][93] = 5'b01111; w[192][94] = 5'b01111; w[192][95] = 5'b01111; w[192][96] = 5'b01111; w[192][97] = 5'b01111; w[192][98] = 5'b01111; w[192][99] = 5'b01111; w[192][100] = 5'b01111; w[192][101] = 5'b00000; w[192][102] = 5'b01111; w[192][103] = 5'b01111; w[192][104] = 5'b10000; w[192][105] = 5'b10000; w[192][106] = 5'b01111; w[192][107] = 5'b00000; w[192][108] = 5'b00000; w[192][109] = 5'b01111; w[192][110] = 5'b01111; w[192][111] = 5'b01111; w[192][112] = 5'b01111; w[192][113] = 5'b01111; w[192][114] = 5'b01111; w[192][115] = 5'b00000; w[192][116] = 5'b01111; w[192][117] = 5'b01111; w[192][118] = 5'b10000; w[192][119] = 5'b10000; w[192][120] = 5'b00000; w[192][121] = 5'b00000; w[192][122] = 5'b00000; w[192][123] = 5'b01111; w[192][124] = 5'b01111; w[192][125] = 5'b01111; w[192][126] = 5'b01111; w[192][127] = 5'b01111; w[192][128] = 5'b01111; w[192][129] = 5'b00000; w[192][130] = 5'b01111; w[192][131] = 5'b01111; w[192][132] = 5'b00000; w[192][133] = 5'b10000; w[192][134] = 5'b01111; w[192][135] = 5'b01111; w[192][136] = 5'b00000; w[192][137] = 5'b01111; w[192][138] = 5'b01111; w[192][139] = 5'b01111; w[192][140] = 5'b01111; w[192][141] = 5'b01111; w[192][142] = 5'b01111; w[192][143] = 5'b00000; w[192][144] = 5'b00000; w[192][145] = 5'b01111; w[192][146] = 5'b00000; w[192][147] = 5'b10000; w[192][148] = 5'b01111; w[192][149] = 5'b00000; w[192][150] = 5'b00000; w[192][151] = 5'b01111; w[192][152] = 5'b01111; w[192][153] = 5'b01111; w[192][154] = 5'b01111; w[192][155] = 5'b01111; w[192][156] = 5'b01111; w[192][157] = 5'b00000; w[192][158] = 5'b00000; w[192][159] = 5'b00000; w[192][160] = 5'b10000; w[192][161] = 5'b10000; w[192][162] = 5'b10000; w[192][163] = 5'b00000; w[192][164] = 5'b00000; w[192][165] = 5'b01111; w[192][166] = 5'b01111; w[192][167] = 5'b01111; w[192][168] = 5'b01111; w[192][169] = 5'b01111; w[192][170] = 5'b01111; w[192][171] = 5'b01111; w[192][172] = 5'b00000; w[192][173] = 5'b00000; w[192][174] = 5'b10000; w[192][175] = 5'b10000; w[192][176] = 5'b10000; w[192][177] = 5'b00000; w[192][178] = 5'b01111; w[192][179] = 5'b01111; w[192][180] = 5'b01111; w[192][181] = 5'b01111; w[192][182] = 5'b01111; w[192][183] = 5'b01111; w[192][184] = 5'b01111; w[192][185] = 5'b01111; w[192][186] = 5'b01111; w[192][187] = 5'b01111; w[192][188] = 5'b01111; w[192][189] = 5'b01111; w[192][190] = 5'b01111; w[192][191] = 5'b01111; w[192][192] = 5'b00000; w[192][193] = 5'b01111; w[192][194] = 5'b01111; w[192][195] = 5'b01111; w[192][196] = 5'b01111; w[192][197] = 5'b01111; w[192][198] = 5'b01111; w[192][199] = 5'b01111; w[192][200] = 5'b01111; w[192][201] = 5'b01111; w[192][202] = 5'b01111; w[192][203] = 5'b01111; w[192][204] = 5'b01111; w[192][205] = 5'b01111; w[192][206] = 5'b01111; w[192][207] = 5'b01111; w[192][208] = 5'b01111; w[192][209] = 5'b01111; 
w[193][0] = 5'b01111; w[193][1] = 5'b01111; w[193][2] = 5'b01111; w[193][3] = 5'b01111; w[193][4] = 5'b01111; w[193][5] = 5'b01111; w[193][6] = 5'b01111; w[193][7] = 5'b01111; w[193][8] = 5'b01111; w[193][9] = 5'b01111; w[193][10] = 5'b01111; w[193][11] = 5'b01111; w[193][12] = 5'b01111; w[193][13] = 5'b01111; w[193][14] = 5'b01111; w[193][15] = 5'b01111; w[193][16] = 5'b01111; w[193][17] = 5'b01111; w[193][18] = 5'b01111; w[193][19] = 5'b01111; w[193][20] = 5'b01111; w[193][21] = 5'b01111; w[193][22] = 5'b01111; w[193][23] = 5'b01111; w[193][24] = 5'b01111; w[193][25] = 5'b01111; w[193][26] = 5'b01111; w[193][27] = 5'b01111; w[193][28] = 5'b01111; w[193][29] = 5'b01111; w[193][30] = 5'b01111; w[193][31] = 5'b00000; w[193][32] = 5'b10000; w[193][33] = 5'b10000; w[193][34] = 5'b10000; w[193][35] = 5'b10000; w[193][36] = 5'b10000; w[193][37] = 5'b10000; w[193][38] = 5'b00000; w[193][39] = 5'b01111; w[193][40] = 5'b01111; w[193][41] = 5'b01111; w[193][42] = 5'b01111; w[193][43] = 5'b01111; w[193][44] = 5'b01111; w[193][45] = 5'b10000; w[193][46] = 5'b10000; w[193][47] = 5'b10000; w[193][48] = 5'b10000; w[193][49] = 5'b10000; w[193][50] = 5'b10000; w[193][51] = 5'b10000; w[193][52] = 5'b10000; w[193][53] = 5'b01111; w[193][54] = 5'b01111; w[193][55] = 5'b01111; w[193][56] = 5'b01111; w[193][57] = 5'b01111; w[193][58] = 5'b01111; w[193][59] = 5'b00000; w[193][60] = 5'b00000; w[193][61] = 5'b01111; w[193][62] = 5'b10000; w[193][63] = 5'b00000; w[193][64] = 5'b01111; w[193][65] = 5'b00000; w[193][66] = 5'b00000; w[193][67] = 5'b01111; w[193][68] = 5'b01111; w[193][69] = 5'b01111; w[193][70] = 5'b01111; w[193][71] = 5'b01111; w[193][72] = 5'b01111; w[193][73] = 5'b00000; w[193][74] = 5'b01111; w[193][75] = 5'b01111; w[193][76] = 5'b10000; w[193][77] = 5'b00000; w[193][78] = 5'b01111; w[193][79] = 5'b01111; w[193][80] = 5'b00000; w[193][81] = 5'b01111; w[193][82] = 5'b01111; w[193][83] = 5'b01111; w[193][84] = 5'b01111; w[193][85] = 5'b01111; w[193][86] = 5'b01111; w[193][87] = 5'b00000; w[193][88] = 5'b01111; w[193][89] = 5'b01111; w[193][90] = 5'b10000; w[193][91] = 5'b10000; w[193][92] = 5'b01111; w[193][93] = 5'b01111; w[193][94] = 5'b01111; w[193][95] = 5'b01111; w[193][96] = 5'b01111; w[193][97] = 5'b01111; w[193][98] = 5'b01111; w[193][99] = 5'b01111; w[193][100] = 5'b01111; w[193][101] = 5'b00000; w[193][102] = 5'b01111; w[193][103] = 5'b01111; w[193][104] = 5'b10000; w[193][105] = 5'b10000; w[193][106] = 5'b01111; w[193][107] = 5'b00000; w[193][108] = 5'b00000; w[193][109] = 5'b01111; w[193][110] = 5'b01111; w[193][111] = 5'b01111; w[193][112] = 5'b01111; w[193][113] = 5'b01111; w[193][114] = 5'b01111; w[193][115] = 5'b00000; w[193][116] = 5'b01111; w[193][117] = 5'b01111; w[193][118] = 5'b10000; w[193][119] = 5'b10000; w[193][120] = 5'b00000; w[193][121] = 5'b00000; w[193][122] = 5'b00000; w[193][123] = 5'b01111; w[193][124] = 5'b01111; w[193][125] = 5'b01111; w[193][126] = 5'b01111; w[193][127] = 5'b01111; w[193][128] = 5'b01111; w[193][129] = 5'b00000; w[193][130] = 5'b01111; w[193][131] = 5'b01111; w[193][132] = 5'b00000; w[193][133] = 5'b10000; w[193][134] = 5'b01111; w[193][135] = 5'b01111; w[193][136] = 5'b00000; w[193][137] = 5'b01111; w[193][138] = 5'b01111; w[193][139] = 5'b01111; w[193][140] = 5'b01111; w[193][141] = 5'b01111; w[193][142] = 5'b01111; w[193][143] = 5'b00000; w[193][144] = 5'b00000; w[193][145] = 5'b01111; w[193][146] = 5'b00000; w[193][147] = 5'b10000; w[193][148] = 5'b01111; w[193][149] = 5'b00000; w[193][150] = 5'b00000; w[193][151] = 5'b01111; w[193][152] = 5'b01111; w[193][153] = 5'b01111; w[193][154] = 5'b01111; w[193][155] = 5'b01111; w[193][156] = 5'b01111; w[193][157] = 5'b00000; w[193][158] = 5'b00000; w[193][159] = 5'b00000; w[193][160] = 5'b10000; w[193][161] = 5'b10000; w[193][162] = 5'b10000; w[193][163] = 5'b00000; w[193][164] = 5'b00000; w[193][165] = 5'b01111; w[193][166] = 5'b01111; w[193][167] = 5'b01111; w[193][168] = 5'b01111; w[193][169] = 5'b01111; w[193][170] = 5'b01111; w[193][171] = 5'b01111; w[193][172] = 5'b00000; w[193][173] = 5'b00000; w[193][174] = 5'b10000; w[193][175] = 5'b10000; w[193][176] = 5'b10000; w[193][177] = 5'b00000; w[193][178] = 5'b01111; w[193][179] = 5'b01111; w[193][180] = 5'b01111; w[193][181] = 5'b01111; w[193][182] = 5'b01111; w[193][183] = 5'b01111; w[193][184] = 5'b01111; w[193][185] = 5'b01111; w[193][186] = 5'b01111; w[193][187] = 5'b01111; w[193][188] = 5'b01111; w[193][189] = 5'b01111; w[193][190] = 5'b01111; w[193][191] = 5'b01111; w[193][192] = 5'b01111; w[193][193] = 5'b00000; w[193][194] = 5'b01111; w[193][195] = 5'b01111; w[193][196] = 5'b01111; w[193][197] = 5'b01111; w[193][198] = 5'b01111; w[193][199] = 5'b01111; w[193][200] = 5'b01111; w[193][201] = 5'b01111; w[193][202] = 5'b01111; w[193][203] = 5'b01111; w[193][204] = 5'b01111; w[193][205] = 5'b01111; w[193][206] = 5'b01111; w[193][207] = 5'b01111; w[193][208] = 5'b01111; w[193][209] = 5'b01111; 
w[194][0] = 5'b01111; w[194][1] = 5'b01111; w[194][2] = 5'b01111; w[194][3] = 5'b01111; w[194][4] = 5'b01111; w[194][5] = 5'b01111; w[194][6] = 5'b01111; w[194][7] = 5'b01111; w[194][8] = 5'b01111; w[194][9] = 5'b01111; w[194][10] = 5'b01111; w[194][11] = 5'b01111; w[194][12] = 5'b01111; w[194][13] = 5'b01111; w[194][14] = 5'b01111; w[194][15] = 5'b01111; w[194][16] = 5'b01111; w[194][17] = 5'b01111; w[194][18] = 5'b01111; w[194][19] = 5'b01111; w[194][20] = 5'b01111; w[194][21] = 5'b01111; w[194][22] = 5'b01111; w[194][23] = 5'b01111; w[194][24] = 5'b01111; w[194][25] = 5'b01111; w[194][26] = 5'b01111; w[194][27] = 5'b01111; w[194][28] = 5'b01111; w[194][29] = 5'b01111; w[194][30] = 5'b01111; w[194][31] = 5'b00000; w[194][32] = 5'b10000; w[194][33] = 5'b10000; w[194][34] = 5'b10000; w[194][35] = 5'b10000; w[194][36] = 5'b10000; w[194][37] = 5'b10000; w[194][38] = 5'b00000; w[194][39] = 5'b01111; w[194][40] = 5'b01111; w[194][41] = 5'b01111; w[194][42] = 5'b01111; w[194][43] = 5'b01111; w[194][44] = 5'b01111; w[194][45] = 5'b10000; w[194][46] = 5'b10000; w[194][47] = 5'b10000; w[194][48] = 5'b10000; w[194][49] = 5'b10000; w[194][50] = 5'b10000; w[194][51] = 5'b10000; w[194][52] = 5'b10000; w[194][53] = 5'b01111; w[194][54] = 5'b01111; w[194][55] = 5'b01111; w[194][56] = 5'b01111; w[194][57] = 5'b01111; w[194][58] = 5'b01111; w[194][59] = 5'b00000; w[194][60] = 5'b00000; w[194][61] = 5'b01111; w[194][62] = 5'b10000; w[194][63] = 5'b00000; w[194][64] = 5'b01111; w[194][65] = 5'b00000; w[194][66] = 5'b00000; w[194][67] = 5'b01111; w[194][68] = 5'b01111; w[194][69] = 5'b01111; w[194][70] = 5'b01111; w[194][71] = 5'b01111; w[194][72] = 5'b01111; w[194][73] = 5'b00000; w[194][74] = 5'b01111; w[194][75] = 5'b01111; w[194][76] = 5'b10000; w[194][77] = 5'b00000; w[194][78] = 5'b01111; w[194][79] = 5'b01111; w[194][80] = 5'b00000; w[194][81] = 5'b01111; w[194][82] = 5'b01111; w[194][83] = 5'b01111; w[194][84] = 5'b01111; w[194][85] = 5'b01111; w[194][86] = 5'b01111; w[194][87] = 5'b00000; w[194][88] = 5'b01111; w[194][89] = 5'b01111; w[194][90] = 5'b10000; w[194][91] = 5'b10000; w[194][92] = 5'b01111; w[194][93] = 5'b01111; w[194][94] = 5'b01111; w[194][95] = 5'b01111; w[194][96] = 5'b01111; w[194][97] = 5'b01111; w[194][98] = 5'b01111; w[194][99] = 5'b01111; w[194][100] = 5'b01111; w[194][101] = 5'b00000; w[194][102] = 5'b01111; w[194][103] = 5'b01111; w[194][104] = 5'b10000; w[194][105] = 5'b10000; w[194][106] = 5'b01111; w[194][107] = 5'b00000; w[194][108] = 5'b00000; w[194][109] = 5'b01111; w[194][110] = 5'b01111; w[194][111] = 5'b01111; w[194][112] = 5'b01111; w[194][113] = 5'b01111; w[194][114] = 5'b01111; w[194][115] = 5'b00000; w[194][116] = 5'b01111; w[194][117] = 5'b01111; w[194][118] = 5'b10000; w[194][119] = 5'b10000; w[194][120] = 5'b00000; w[194][121] = 5'b00000; w[194][122] = 5'b00000; w[194][123] = 5'b01111; w[194][124] = 5'b01111; w[194][125] = 5'b01111; w[194][126] = 5'b01111; w[194][127] = 5'b01111; w[194][128] = 5'b01111; w[194][129] = 5'b00000; w[194][130] = 5'b01111; w[194][131] = 5'b01111; w[194][132] = 5'b00000; w[194][133] = 5'b10000; w[194][134] = 5'b01111; w[194][135] = 5'b01111; w[194][136] = 5'b00000; w[194][137] = 5'b01111; w[194][138] = 5'b01111; w[194][139] = 5'b01111; w[194][140] = 5'b01111; w[194][141] = 5'b01111; w[194][142] = 5'b01111; w[194][143] = 5'b00000; w[194][144] = 5'b00000; w[194][145] = 5'b01111; w[194][146] = 5'b00000; w[194][147] = 5'b10000; w[194][148] = 5'b01111; w[194][149] = 5'b00000; w[194][150] = 5'b00000; w[194][151] = 5'b01111; w[194][152] = 5'b01111; w[194][153] = 5'b01111; w[194][154] = 5'b01111; w[194][155] = 5'b01111; w[194][156] = 5'b01111; w[194][157] = 5'b00000; w[194][158] = 5'b00000; w[194][159] = 5'b00000; w[194][160] = 5'b10000; w[194][161] = 5'b10000; w[194][162] = 5'b10000; w[194][163] = 5'b00000; w[194][164] = 5'b00000; w[194][165] = 5'b01111; w[194][166] = 5'b01111; w[194][167] = 5'b01111; w[194][168] = 5'b01111; w[194][169] = 5'b01111; w[194][170] = 5'b01111; w[194][171] = 5'b01111; w[194][172] = 5'b00000; w[194][173] = 5'b00000; w[194][174] = 5'b10000; w[194][175] = 5'b10000; w[194][176] = 5'b10000; w[194][177] = 5'b00000; w[194][178] = 5'b01111; w[194][179] = 5'b01111; w[194][180] = 5'b01111; w[194][181] = 5'b01111; w[194][182] = 5'b01111; w[194][183] = 5'b01111; w[194][184] = 5'b01111; w[194][185] = 5'b01111; w[194][186] = 5'b01111; w[194][187] = 5'b01111; w[194][188] = 5'b01111; w[194][189] = 5'b01111; w[194][190] = 5'b01111; w[194][191] = 5'b01111; w[194][192] = 5'b01111; w[194][193] = 5'b01111; w[194][194] = 5'b00000; w[194][195] = 5'b01111; w[194][196] = 5'b01111; w[194][197] = 5'b01111; w[194][198] = 5'b01111; w[194][199] = 5'b01111; w[194][200] = 5'b01111; w[194][201] = 5'b01111; w[194][202] = 5'b01111; w[194][203] = 5'b01111; w[194][204] = 5'b01111; w[194][205] = 5'b01111; w[194][206] = 5'b01111; w[194][207] = 5'b01111; w[194][208] = 5'b01111; w[194][209] = 5'b01111; 
w[195][0] = 5'b01111; w[195][1] = 5'b01111; w[195][2] = 5'b01111; w[195][3] = 5'b01111; w[195][4] = 5'b01111; w[195][5] = 5'b01111; w[195][6] = 5'b01111; w[195][7] = 5'b01111; w[195][8] = 5'b01111; w[195][9] = 5'b01111; w[195][10] = 5'b01111; w[195][11] = 5'b01111; w[195][12] = 5'b01111; w[195][13] = 5'b01111; w[195][14] = 5'b01111; w[195][15] = 5'b01111; w[195][16] = 5'b01111; w[195][17] = 5'b01111; w[195][18] = 5'b01111; w[195][19] = 5'b01111; w[195][20] = 5'b01111; w[195][21] = 5'b01111; w[195][22] = 5'b01111; w[195][23] = 5'b01111; w[195][24] = 5'b01111; w[195][25] = 5'b01111; w[195][26] = 5'b01111; w[195][27] = 5'b01111; w[195][28] = 5'b01111; w[195][29] = 5'b01111; w[195][30] = 5'b01111; w[195][31] = 5'b00000; w[195][32] = 5'b10000; w[195][33] = 5'b10000; w[195][34] = 5'b10000; w[195][35] = 5'b10000; w[195][36] = 5'b10000; w[195][37] = 5'b10000; w[195][38] = 5'b00000; w[195][39] = 5'b01111; w[195][40] = 5'b01111; w[195][41] = 5'b01111; w[195][42] = 5'b01111; w[195][43] = 5'b01111; w[195][44] = 5'b01111; w[195][45] = 5'b10000; w[195][46] = 5'b10000; w[195][47] = 5'b10000; w[195][48] = 5'b10000; w[195][49] = 5'b10000; w[195][50] = 5'b10000; w[195][51] = 5'b10000; w[195][52] = 5'b10000; w[195][53] = 5'b01111; w[195][54] = 5'b01111; w[195][55] = 5'b01111; w[195][56] = 5'b01111; w[195][57] = 5'b01111; w[195][58] = 5'b01111; w[195][59] = 5'b00000; w[195][60] = 5'b00000; w[195][61] = 5'b01111; w[195][62] = 5'b10000; w[195][63] = 5'b00000; w[195][64] = 5'b01111; w[195][65] = 5'b00000; w[195][66] = 5'b00000; w[195][67] = 5'b01111; w[195][68] = 5'b01111; w[195][69] = 5'b01111; w[195][70] = 5'b01111; w[195][71] = 5'b01111; w[195][72] = 5'b01111; w[195][73] = 5'b00000; w[195][74] = 5'b01111; w[195][75] = 5'b01111; w[195][76] = 5'b10000; w[195][77] = 5'b00000; w[195][78] = 5'b01111; w[195][79] = 5'b01111; w[195][80] = 5'b00000; w[195][81] = 5'b01111; w[195][82] = 5'b01111; w[195][83] = 5'b01111; w[195][84] = 5'b01111; w[195][85] = 5'b01111; w[195][86] = 5'b01111; w[195][87] = 5'b00000; w[195][88] = 5'b01111; w[195][89] = 5'b01111; w[195][90] = 5'b10000; w[195][91] = 5'b10000; w[195][92] = 5'b01111; w[195][93] = 5'b01111; w[195][94] = 5'b01111; w[195][95] = 5'b01111; w[195][96] = 5'b01111; w[195][97] = 5'b01111; w[195][98] = 5'b01111; w[195][99] = 5'b01111; w[195][100] = 5'b01111; w[195][101] = 5'b00000; w[195][102] = 5'b01111; w[195][103] = 5'b01111; w[195][104] = 5'b10000; w[195][105] = 5'b10000; w[195][106] = 5'b01111; w[195][107] = 5'b00000; w[195][108] = 5'b00000; w[195][109] = 5'b01111; w[195][110] = 5'b01111; w[195][111] = 5'b01111; w[195][112] = 5'b01111; w[195][113] = 5'b01111; w[195][114] = 5'b01111; w[195][115] = 5'b00000; w[195][116] = 5'b01111; w[195][117] = 5'b01111; w[195][118] = 5'b10000; w[195][119] = 5'b10000; w[195][120] = 5'b00000; w[195][121] = 5'b00000; w[195][122] = 5'b00000; w[195][123] = 5'b01111; w[195][124] = 5'b01111; w[195][125] = 5'b01111; w[195][126] = 5'b01111; w[195][127] = 5'b01111; w[195][128] = 5'b01111; w[195][129] = 5'b00000; w[195][130] = 5'b01111; w[195][131] = 5'b01111; w[195][132] = 5'b00000; w[195][133] = 5'b10000; w[195][134] = 5'b01111; w[195][135] = 5'b01111; w[195][136] = 5'b00000; w[195][137] = 5'b01111; w[195][138] = 5'b01111; w[195][139] = 5'b01111; w[195][140] = 5'b01111; w[195][141] = 5'b01111; w[195][142] = 5'b01111; w[195][143] = 5'b00000; w[195][144] = 5'b00000; w[195][145] = 5'b01111; w[195][146] = 5'b00000; w[195][147] = 5'b10000; w[195][148] = 5'b01111; w[195][149] = 5'b00000; w[195][150] = 5'b00000; w[195][151] = 5'b01111; w[195][152] = 5'b01111; w[195][153] = 5'b01111; w[195][154] = 5'b01111; w[195][155] = 5'b01111; w[195][156] = 5'b01111; w[195][157] = 5'b00000; w[195][158] = 5'b00000; w[195][159] = 5'b00000; w[195][160] = 5'b10000; w[195][161] = 5'b10000; w[195][162] = 5'b10000; w[195][163] = 5'b00000; w[195][164] = 5'b00000; w[195][165] = 5'b01111; w[195][166] = 5'b01111; w[195][167] = 5'b01111; w[195][168] = 5'b01111; w[195][169] = 5'b01111; w[195][170] = 5'b01111; w[195][171] = 5'b01111; w[195][172] = 5'b00000; w[195][173] = 5'b00000; w[195][174] = 5'b10000; w[195][175] = 5'b10000; w[195][176] = 5'b10000; w[195][177] = 5'b00000; w[195][178] = 5'b01111; w[195][179] = 5'b01111; w[195][180] = 5'b01111; w[195][181] = 5'b01111; w[195][182] = 5'b01111; w[195][183] = 5'b01111; w[195][184] = 5'b01111; w[195][185] = 5'b01111; w[195][186] = 5'b01111; w[195][187] = 5'b01111; w[195][188] = 5'b01111; w[195][189] = 5'b01111; w[195][190] = 5'b01111; w[195][191] = 5'b01111; w[195][192] = 5'b01111; w[195][193] = 5'b01111; w[195][194] = 5'b01111; w[195][195] = 5'b00000; w[195][196] = 5'b01111; w[195][197] = 5'b01111; w[195][198] = 5'b01111; w[195][199] = 5'b01111; w[195][200] = 5'b01111; w[195][201] = 5'b01111; w[195][202] = 5'b01111; w[195][203] = 5'b01111; w[195][204] = 5'b01111; w[195][205] = 5'b01111; w[195][206] = 5'b01111; w[195][207] = 5'b01111; w[195][208] = 5'b01111; w[195][209] = 5'b01111; 
w[196][0] = 5'b01111; w[196][1] = 5'b01111; w[196][2] = 5'b01111; w[196][3] = 5'b01111; w[196][4] = 5'b01111; w[196][5] = 5'b01111; w[196][6] = 5'b01111; w[196][7] = 5'b01111; w[196][8] = 5'b01111; w[196][9] = 5'b01111; w[196][10] = 5'b01111; w[196][11] = 5'b01111; w[196][12] = 5'b01111; w[196][13] = 5'b01111; w[196][14] = 5'b01111; w[196][15] = 5'b01111; w[196][16] = 5'b01111; w[196][17] = 5'b01111; w[196][18] = 5'b01111; w[196][19] = 5'b01111; w[196][20] = 5'b01111; w[196][21] = 5'b01111; w[196][22] = 5'b01111; w[196][23] = 5'b01111; w[196][24] = 5'b01111; w[196][25] = 5'b01111; w[196][26] = 5'b01111; w[196][27] = 5'b01111; w[196][28] = 5'b01111; w[196][29] = 5'b01111; w[196][30] = 5'b01111; w[196][31] = 5'b00000; w[196][32] = 5'b10000; w[196][33] = 5'b10000; w[196][34] = 5'b10000; w[196][35] = 5'b10000; w[196][36] = 5'b10000; w[196][37] = 5'b10000; w[196][38] = 5'b00000; w[196][39] = 5'b01111; w[196][40] = 5'b01111; w[196][41] = 5'b01111; w[196][42] = 5'b01111; w[196][43] = 5'b01111; w[196][44] = 5'b01111; w[196][45] = 5'b10000; w[196][46] = 5'b10000; w[196][47] = 5'b10000; w[196][48] = 5'b10000; w[196][49] = 5'b10000; w[196][50] = 5'b10000; w[196][51] = 5'b10000; w[196][52] = 5'b10000; w[196][53] = 5'b01111; w[196][54] = 5'b01111; w[196][55] = 5'b01111; w[196][56] = 5'b01111; w[196][57] = 5'b01111; w[196][58] = 5'b01111; w[196][59] = 5'b00000; w[196][60] = 5'b00000; w[196][61] = 5'b01111; w[196][62] = 5'b10000; w[196][63] = 5'b00000; w[196][64] = 5'b01111; w[196][65] = 5'b00000; w[196][66] = 5'b00000; w[196][67] = 5'b01111; w[196][68] = 5'b01111; w[196][69] = 5'b01111; w[196][70] = 5'b01111; w[196][71] = 5'b01111; w[196][72] = 5'b01111; w[196][73] = 5'b00000; w[196][74] = 5'b01111; w[196][75] = 5'b01111; w[196][76] = 5'b10000; w[196][77] = 5'b00000; w[196][78] = 5'b01111; w[196][79] = 5'b01111; w[196][80] = 5'b00000; w[196][81] = 5'b01111; w[196][82] = 5'b01111; w[196][83] = 5'b01111; w[196][84] = 5'b01111; w[196][85] = 5'b01111; w[196][86] = 5'b01111; w[196][87] = 5'b00000; w[196][88] = 5'b01111; w[196][89] = 5'b01111; w[196][90] = 5'b10000; w[196][91] = 5'b10000; w[196][92] = 5'b01111; w[196][93] = 5'b01111; w[196][94] = 5'b01111; w[196][95] = 5'b01111; w[196][96] = 5'b01111; w[196][97] = 5'b01111; w[196][98] = 5'b01111; w[196][99] = 5'b01111; w[196][100] = 5'b01111; w[196][101] = 5'b00000; w[196][102] = 5'b01111; w[196][103] = 5'b01111; w[196][104] = 5'b10000; w[196][105] = 5'b10000; w[196][106] = 5'b01111; w[196][107] = 5'b00000; w[196][108] = 5'b00000; w[196][109] = 5'b01111; w[196][110] = 5'b01111; w[196][111] = 5'b01111; w[196][112] = 5'b01111; w[196][113] = 5'b01111; w[196][114] = 5'b01111; w[196][115] = 5'b00000; w[196][116] = 5'b01111; w[196][117] = 5'b01111; w[196][118] = 5'b10000; w[196][119] = 5'b10000; w[196][120] = 5'b00000; w[196][121] = 5'b00000; w[196][122] = 5'b00000; w[196][123] = 5'b01111; w[196][124] = 5'b01111; w[196][125] = 5'b01111; w[196][126] = 5'b01111; w[196][127] = 5'b01111; w[196][128] = 5'b01111; w[196][129] = 5'b00000; w[196][130] = 5'b01111; w[196][131] = 5'b01111; w[196][132] = 5'b00000; w[196][133] = 5'b10000; w[196][134] = 5'b01111; w[196][135] = 5'b01111; w[196][136] = 5'b00000; w[196][137] = 5'b01111; w[196][138] = 5'b01111; w[196][139] = 5'b01111; w[196][140] = 5'b01111; w[196][141] = 5'b01111; w[196][142] = 5'b01111; w[196][143] = 5'b00000; w[196][144] = 5'b00000; w[196][145] = 5'b01111; w[196][146] = 5'b00000; w[196][147] = 5'b10000; w[196][148] = 5'b01111; w[196][149] = 5'b00000; w[196][150] = 5'b00000; w[196][151] = 5'b01111; w[196][152] = 5'b01111; w[196][153] = 5'b01111; w[196][154] = 5'b01111; w[196][155] = 5'b01111; w[196][156] = 5'b01111; w[196][157] = 5'b00000; w[196][158] = 5'b00000; w[196][159] = 5'b00000; w[196][160] = 5'b10000; w[196][161] = 5'b10000; w[196][162] = 5'b10000; w[196][163] = 5'b00000; w[196][164] = 5'b00000; w[196][165] = 5'b01111; w[196][166] = 5'b01111; w[196][167] = 5'b01111; w[196][168] = 5'b01111; w[196][169] = 5'b01111; w[196][170] = 5'b01111; w[196][171] = 5'b01111; w[196][172] = 5'b00000; w[196][173] = 5'b00000; w[196][174] = 5'b10000; w[196][175] = 5'b10000; w[196][176] = 5'b10000; w[196][177] = 5'b00000; w[196][178] = 5'b01111; w[196][179] = 5'b01111; w[196][180] = 5'b01111; w[196][181] = 5'b01111; w[196][182] = 5'b01111; w[196][183] = 5'b01111; w[196][184] = 5'b01111; w[196][185] = 5'b01111; w[196][186] = 5'b01111; w[196][187] = 5'b01111; w[196][188] = 5'b01111; w[196][189] = 5'b01111; w[196][190] = 5'b01111; w[196][191] = 5'b01111; w[196][192] = 5'b01111; w[196][193] = 5'b01111; w[196][194] = 5'b01111; w[196][195] = 5'b01111; w[196][196] = 5'b00000; w[196][197] = 5'b01111; w[196][198] = 5'b01111; w[196][199] = 5'b01111; w[196][200] = 5'b01111; w[196][201] = 5'b01111; w[196][202] = 5'b01111; w[196][203] = 5'b01111; w[196][204] = 5'b01111; w[196][205] = 5'b01111; w[196][206] = 5'b01111; w[196][207] = 5'b01111; w[196][208] = 5'b01111; w[196][209] = 5'b01111; 
w[197][0] = 5'b01111; w[197][1] = 5'b01111; w[197][2] = 5'b01111; w[197][3] = 5'b01111; w[197][4] = 5'b01111; w[197][5] = 5'b01111; w[197][6] = 5'b01111; w[197][7] = 5'b01111; w[197][8] = 5'b01111; w[197][9] = 5'b01111; w[197][10] = 5'b01111; w[197][11] = 5'b01111; w[197][12] = 5'b01111; w[197][13] = 5'b01111; w[197][14] = 5'b01111; w[197][15] = 5'b01111; w[197][16] = 5'b01111; w[197][17] = 5'b01111; w[197][18] = 5'b01111; w[197][19] = 5'b01111; w[197][20] = 5'b01111; w[197][21] = 5'b01111; w[197][22] = 5'b01111; w[197][23] = 5'b01111; w[197][24] = 5'b01111; w[197][25] = 5'b01111; w[197][26] = 5'b01111; w[197][27] = 5'b01111; w[197][28] = 5'b01111; w[197][29] = 5'b01111; w[197][30] = 5'b01111; w[197][31] = 5'b00000; w[197][32] = 5'b10000; w[197][33] = 5'b10000; w[197][34] = 5'b10000; w[197][35] = 5'b10000; w[197][36] = 5'b10000; w[197][37] = 5'b10000; w[197][38] = 5'b00000; w[197][39] = 5'b01111; w[197][40] = 5'b01111; w[197][41] = 5'b01111; w[197][42] = 5'b01111; w[197][43] = 5'b01111; w[197][44] = 5'b01111; w[197][45] = 5'b10000; w[197][46] = 5'b10000; w[197][47] = 5'b10000; w[197][48] = 5'b10000; w[197][49] = 5'b10000; w[197][50] = 5'b10000; w[197][51] = 5'b10000; w[197][52] = 5'b10000; w[197][53] = 5'b01111; w[197][54] = 5'b01111; w[197][55] = 5'b01111; w[197][56] = 5'b01111; w[197][57] = 5'b01111; w[197][58] = 5'b01111; w[197][59] = 5'b00000; w[197][60] = 5'b00000; w[197][61] = 5'b01111; w[197][62] = 5'b10000; w[197][63] = 5'b00000; w[197][64] = 5'b01111; w[197][65] = 5'b00000; w[197][66] = 5'b00000; w[197][67] = 5'b01111; w[197][68] = 5'b01111; w[197][69] = 5'b01111; w[197][70] = 5'b01111; w[197][71] = 5'b01111; w[197][72] = 5'b01111; w[197][73] = 5'b00000; w[197][74] = 5'b01111; w[197][75] = 5'b01111; w[197][76] = 5'b10000; w[197][77] = 5'b00000; w[197][78] = 5'b01111; w[197][79] = 5'b01111; w[197][80] = 5'b00000; w[197][81] = 5'b01111; w[197][82] = 5'b01111; w[197][83] = 5'b01111; w[197][84] = 5'b01111; w[197][85] = 5'b01111; w[197][86] = 5'b01111; w[197][87] = 5'b00000; w[197][88] = 5'b01111; w[197][89] = 5'b01111; w[197][90] = 5'b10000; w[197][91] = 5'b10000; w[197][92] = 5'b01111; w[197][93] = 5'b01111; w[197][94] = 5'b01111; w[197][95] = 5'b01111; w[197][96] = 5'b01111; w[197][97] = 5'b01111; w[197][98] = 5'b01111; w[197][99] = 5'b01111; w[197][100] = 5'b01111; w[197][101] = 5'b00000; w[197][102] = 5'b01111; w[197][103] = 5'b01111; w[197][104] = 5'b10000; w[197][105] = 5'b10000; w[197][106] = 5'b01111; w[197][107] = 5'b00000; w[197][108] = 5'b00000; w[197][109] = 5'b01111; w[197][110] = 5'b01111; w[197][111] = 5'b01111; w[197][112] = 5'b01111; w[197][113] = 5'b01111; w[197][114] = 5'b01111; w[197][115] = 5'b00000; w[197][116] = 5'b01111; w[197][117] = 5'b01111; w[197][118] = 5'b10000; w[197][119] = 5'b10000; w[197][120] = 5'b00000; w[197][121] = 5'b00000; w[197][122] = 5'b00000; w[197][123] = 5'b01111; w[197][124] = 5'b01111; w[197][125] = 5'b01111; w[197][126] = 5'b01111; w[197][127] = 5'b01111; w[197][128] = 5'b01111; w[197][129] = 5'b00000; w[197][130] = 5'b01111; w[197][131] = 5'b01111; w[197][132] = 5'b00000; w[197][133] = 5'b10000; w[197][134] = 5'b01111; w[197][135] = 5'b01111; w[197][136] = 5'b00000; w[197][137] = 5'b01111; w[197][138] = 5'b01111; w[197][139] = 5'b01111; w[197][140] = 5'b01111; w[197][141] = 5'b01111; w[197][142] = 5'b01111; w[197][143] = 5'b00000; w[197][144] = 5'b00000; w[197][145] = 5'b01111; w[197][146] = 5'b00000; w[197][147] = 5'b10000; w[197][148] = 5'b01111; w[197][149] = 5'b00000; w[197][150] = 5'b00000; w[197][151] = 5'b01111; w[197][152] = 5'b01111; w[197][153] = 5'b01111; w[197][154] = 5'b01111; w[197][155] = 5'b01111; w[197][156] = 5'b01111; w[197][157] = 5'b00000; w[197][158] = 5'b00000; w[197][159] = 5'b00000; w[197][160] = 5'b10000; w[197][161] = 5'b10000; w[197][162] = 5'b10000; w[197][163] = 5'b00000; w[197][164] = 5'b00000; w[197][165] = 5'b01111; w[197][166] = 5'b01111; w[197][167] = 5'b01111; w[197][168] = 5'b01111; w[197][169] = 5'b01111; w[197][170] = 5'b01111; w[197][171] = 5'b01111; w[197][172] = 5'b00000; w[197][173] = 5'b00000; w[197][174] = 5'b10000; w[197][175] = 5'b10000; w[197][176] = 5'b10000; w[197][177] = 5'b00000; w[197][178] = 5'b01111; w[197][179] = 5'b01111; w[197][180] = 5'b01111; w[197][181] = 5'b01111; w[197][182] = 5'b01111; w[197][183] = 5'b01111; w[197][184] = 5'b01111; w[197][185] = 5'b01111; w[197][186] = 5'b01111; w[197][187] = 5'b01111; w[197][188] = 5'b01111; w[197][189] = 5'b01111; w[197][190] = 5'b01111; w[197][191] = 5'b01111; w[197][192] = 5'b01111; w[197][193] = 5'b01111; w[197][194] = 5'b01111; w[197][195] = 5'b01111; w[197][196] = 5'b01111; w[197][197] = 5'b00000; w[197][198] = 5'b01111; w[197][199] = 5'b01111; w[197][200] = 5'b01111; w[197][201] = 5'b01111; w[197][202] = 5'b01111; w[197][203] = 5'b01111; w[197][204] = 5'b01111; w[197][205] = 5'b01111; w[197][206] = 5'b01111; w[197][207] = 5'b01111; w[197][208] = 5'b01111; w[197][209] = 5'b01111; 
w[198][0] = 5'b01111; w[198][1] = 5'b01111; w[198][2] = 5'b01111; w[198][3] = 5'b01111; w[198][4] = 5'b01111; w[198][5] = 5'b01111; w[198][6] = 5'b01111; w[198][7] = 5'b01111; w[198][8] = 5'b01111; w[198][9] = 5'b01111; w[198][10] = 5'b01111; w[198][11] = 5'b01111; w[198][12] = 5'b01111; w[198][13] = 5'b01111; w[198][14] = 5'b01111; w[198][15] = 5'b01111; w[198][16] = 5'b01111; w[198][17] = 5'b01111; w[198][18] = 5'b01111; w[198][19] = 5'b01111; w[198][20] = 5'b01111; w[198][21] = 5'b01111; w[198][22] = 5'b01111; w[198][23] = 5'b01111; w[198][24] = 5'b01111; w[198][25] = 5'b01111; w[198][26] = 5'b01111; w[198][27] = 5'b01111; w[198][28] = 5'b01111; w[198][29] = 5'b01111; w[198][30] = 5'b01111; w[198][31] = 5'b00000; w[198][32] = 5'b10000; w[198][33] = 5'b10000; w[198][34] = 5'b10000; w[198][35] = 5'b10000; w[198][36] = 5'b10000; w[198][37] = 5'b10000; w[198][38] = 5'b00000; w[198][39] = 5'b01111; w[198][40] = 5'b01111; w[198][41] = 5'b01111; w[198][42] = 5'b01111; w[198][43] = 5'b01111; w[198][44] = 5'b01111; w[198][45] = 5'b10000; w[198][46] = 5'b10000; w[198][47] = 5'b10000; w[198][48] = 5'b10000; w[198][49] = 5'b10000; w[198][50] = 5'b10000; w[198][51] = 5'b10000; w[198][52] = 5'b10000; w[198][53] = 5'b01111; w[198][54] = 5'b01111; w[198][55] = 5'b01111; w[198][56] = 5'b01111; w[198][57] = 5'b01111; w[198][58] = 5'b01111; w[198][59] = 5'b00000; w[198][60] = 5'b00000; w[198][61] = 5'b01111; w[198][62] = 5'b10000; w[198][63] = 5'b00000; w[198][64] = 5'b01111; w[198][65] = 5'b00000; w[198][66] = 5'b00000; w[198][67] = 5'b01111; w[198][68] = 5'b01111; w[198][69] = 5'b01111; w[198][70] = 5'b01111; w[198][71] = 5'b01111; w[198][72] = 5'b01111; w[198][73] = 5'b00000; w[198][74] = 5'b01111; w[198][75] = 5'b01111; w[198][76] = 5'b10000; w[198][77] = 5'b00000; w[198][78] = 5'b01111; w[198][79] = 5'b01111; w[198][80] = 5'b00000; w[198][81] = 5'b01111; w[198][82] = 5'b01111; w[198][83] = 5'b01111; w[198][84] = 5'b01111; w[198][85] = 5'b01111; w[198][86] = 5'b01111; w[198][87] = 5'b00000; w[198][88] = 5'b01111; w[198][89] = 5'b01111; w[198][90] = 5'b10000; w[198][91] = 5'b10000; w[198][92] = 5'b01111; w[198][93] = 5'b01111; w[198][94] = 5'b01111; w[198][95] = 5'b01111; w[198][96] = 5'b01111; w[198][97] = 5'b01111; w[198][98] = 5'b01111; w[198][99] = 5'b01111; w[198][100] = 5'b01111; w[198][101] = 5'b00000; w[198][102] = 5'b01111; w[198][103] = 5'b01111; w[198][104] = 5'b10000; w[198][105] = 5'b10000; w[198][106] = 5'b01111; w[198][107] = 5'b00000; w[198][108] = 5'b00000; w[198][109] = 5'b01111; w[198][110] = 5'b01111; w[198][111] = 5'b01111; w[198][112] = 5'b01111; w[198][113] = 5'b01111; w[198][114] = 5'b01111; w[198][115] = 5'b00000; w[198][116] = 5'b01111; w[198][117] = 5'b01111; w[198][118] = 5'b10000; w[198][119] = 5'b10000; w[198][120] = 5'b00000; w[198][121] = 5'b00000; w[198][122] = 5'b00000; w[198][123] = 5'b01111; w[198][124] = 5'b01111; w[198][125] = 5'b01111; w[198][126] = 5'b01111; w[198][127] = 5'b01111; w[198][128] = 5'b01111; w[198][129] = 5'b00000; w[198][130] = 5'b01111; w[198][131] = 5'b01111; w[198][132] = 5'b00000; w[198][133] = 5'b10000; w[198][134] = 5'b01111; w[198][135] = 5'b01111; w[198][136] = 5'b00000; w[198][137] = 5'b01111; w[198][138] = 5'b01111; w[198][139] = 5'b01111; w[198][140] = 5'b01111; w[198][141] = 5'b01111; w[198][142] = 5'b01111; w[198][143] = 5'b00000; w[198][144] = 5'b00000; w[198][145] = 5'b01111; w[198][146] = 5'b00000; w[198][147] = 5'b10000; w[198][148] = 5'b01111; w[198][149] = 5'b00000; w[198][150] = 5'b00000; w[198][151] = 5'b01111; w[198][152] = 5'b01111; w[198][153] = 5'b01111; w[198][154] = 5'b01111; w[198][155] = 5'b01111; w[198][156] = 5'b01111; w[198][157] = 5'b00000; w[198][158] = 5'b00000; w[198][159] = 5'b00000; w[198][160] = 5'b10000; w[198][161] = 5'b10000; w[198][162] = 5'b10000; w[198][163] = 5'b00000; w[198][164] = 5'b00000; w[198][165] = 5'b01111; w[198][166] = 5'b01111; w[198][167] = 5'b01111; w[198][168] = 5'b01111; w[198][169] = 5'b01111; w[198][170] = 5'b01111; w[198][171] = 5'b01111; w[198][172] = 5'b00000; w[198][173] = 5'b00000; w[198][174] = 5'b10000; w[198][175] = 5'b10000; w[198][176] = 5'b10000; w[198][177] = 5'b00000; w[198][178] = 5'b01111; w[198][179] = 5'b01111; w[198][180] = 5'b01111; w[198][181] = 5'b01111; w[198][182] = 5'b01111; w[198][183] = 5'b01111; w[198][184] = 5'b01111; w[198][185] = 5'b01111; w[198][186] = 5'b01111; w[198][187] = 5'b01111; w[198][188] = 5'b01111; w[198][189] = 5'b01111; w[198][190] = 5'b01111; w[198][191] = 5'b01111; w[198][192] = 5'b01111; w[198][193] = 5'b01111; w[198][194] = 5'b01111; w[198][195] = 5'b01111; w[198][196] = 5'b01111; w[198][197] = 5'b01111; w[198][198] = 5'b00000; w[198][199] = 5'b01111; w[198][200] = 5'b01111; w[198][201] = 5'b01111; w[198][202] = 5'b01111; w[198][203] = 5'b01111; w[198][204] = 5'b01111; w[198][205] = 5'b01111; w[198][206] = 5'b01111; w[198][207] = 5'b01111; w[198][208] = 5'b01111; w[198][209] = 5'b01111; 
w[199][0] = 5'b01111; w[199][1] = 5'b01111; w[199][2] = 5'b01111; w[199][3] = 5'b01111; w[199][4] = 5'b01111; w[199][5] = 5'b01111; w[199][6] = 5'b01111; w[199][7] = 5'b01111; w[199][8] = 5'b01111; w[199][9] = 5'b01111; w[199][10] = 5'b01111; w[199][11] = 5'b01111; w[199][12] = 5'b01111; w[199][13] = 5'b01111; w[199][14] = 5'b01111; w[199][15] = 5'b01111; w[199][16] = 5'b01111; w[199][17] = 5'b01111; w[199][18] = 5'b01111; w[199][19] = 5'b01111; w[199][20] = 5'b01111; w[199][21] = 5'b01111; w[199][22] = 5'b01111; w[199][23] = 5'b01111; w[199][24] = 5'b01111; w[199][25] = 5'b01111; w[199][26] = 5'b01111; w[199][27] = 5'b01111; w[199][28] = 5'b01111; w[199][29] = 5'b01111; w[199][30] = 5'b01111; w[199][31] = 5'b00000; w[199][32] = 5'b10000; w[199][33] = 5'b10000; w[199][34] = 5'b10000; w[199][35] = 5'b10000; w[199][36] = 5'b10000; w[199][37] = 5'b10000; w[199][38] = 5'b00000; w[199][39] = 5'b01111; w[199][40] = 5'b01111; w[199][41] = 5'b01111; w[199][42] = 5'b01111; w[199][43] = 5'b01111; w[199][44] = 5'b01111; w[199][45] = 5'b10000; w[199][46] = 5'b10000; w[199][47] = 5'b10000; w[199][48] = 5'b10000; w[199][49] = 5'b10000; w[199][50] = 5'b10000; w[199][51] = 5'b10000; w[199][52] = 5'b10000; w[199][53] = 5'b01111; w[199][54] = 5'b01111; w[199][55] = 5'b01111; w[199][56] = 5'b01111; w[199][57] = 5'b01111; w[199][58] = 5'b01111; w[199][59] = 5'b00000; w[199][60] = 5'b00000; w[199][61] = 5'b01111; w[199][62] = 5'b10000; w[199][63] = 5'b00000; w[199][64] = 5'b01111; w[199][65] = 5'b00000; w[199][66] = 5'b00000; w[199][67] = 5'b01111; w[199][68] = 5'b01111; w[199][69] = 5'b01111; w[199][70] = 5'b01111; w[199][71] = 5'b01111; w[199][72] = 5'b01111; w[199][73] = 5'b00000; w[199][74] = 5'b01111; w[199][75] = 5'b01111; w[199][76] = 5'b10000; w[199][77] = 5'b00000; w[199][78] = 5'b01111; w[199][79] = 5'b01111; w[199][80] = 5'b00000; w[199][81] = 5'b01111; w[199][82] = 5'b01111; w[199][83] = 5'b01111; w[199][84] = 5'b01111; w[199][85] = 5'b01111; w[199][86] = 5'b01111; w[199][87] = 5'b00000; w[199][88] = 5'b01111; w[199][89] = 5'b01111; w[199][90] = 5'b10000; w[199][91] = 5'b10000; w[199][92] = 5'b01111; w[199][93] = 5'b01111; w[199][94] = 5'b01111; w[199][95] = 5'b01111; w[199][96] = 5'b01111; w[199][97] = 5'b01111; w[199][98] = 5'b01111; w[199][99] = 5'b01111; w[199][100] = 5'b01111; w[199][101] = 5'b00000; w[199][102] = 5'b01111; w[199][103] = 5'b01111; w[199][104] = 5'b10000; w[199][105] = 5'b10000; w[199][106] = 5'b01111; w[199][107] = 5'b00000; w[199][108] = 5'b00000; w[199][109] = 5'b01111; w[199][110] = 5'b01111; w[199][111] = 5'b01111; w[199][112] = 5'b01111; w[199][113] = 5'b01111; w[199][114] = 5'b01111; w[199][115] = 5'b00000; w[199][116] = 5'b01111; w[199][117] = 5'b01111; w[199][118] = 5'b10000; w[199][119] = 5'b10000; w[199][120] = 5'b00000; w[199][121] = 5'b00000; w[199][122] = 5'b00000; w[199][123] = 5'b01111; w[199][124] = 5'b01111; w[199][125] = 5'b01111; w[199][126] = 5'b01111; w[199][127] = 5'b01111; w[199][128] = 5'b01111; w[199][129] = 5'b00000; w[199][130] = 5'b01111; w[199][131] = 5'b01111; w[199][132] = 5'b00000; w[199][133] = 5'b10000; w[199][134] = 5'b01111; w[199][135] = 5'b01111; w[199][136] = 5'b00000; w[199][137] = 5'b01111; w[199][138] = 5'b01111; w[199][139] = 5'b01111; w[199][140] = 5'b01111; w[199][141] = 5'b01111; w[199][142] = 5'b01111; w[199][143] = 5'b00000; w[199][144] = 5'b00000; w[199][145] = 5'b01111; w[199][146] = 5'b00000; w[199][147] = 5'b10000; w[199][148] = 5'b01111; w[199][149] = 5'b00000; w[199][150] = 5'b00000; w[199][151] = 5'b01111; w[199][152] = 5'b01111; w[199][153] = 5'b01111; w[199][154] = 5'b01111; w[199][155] = 5'b01111; w[199][156] = 5'b01111; w[199][157] = 5'b00000; w[199][158] = 5'b00000; w[199][159] = 5'b00000; w[199][160] = 5'b10000; w[199][161] = 5'b10000; w[199][162] = 5'b10000; w[199][163] = 5'b00000; w[199][164] = 5'b00000; w[199][165] = 5'b01111; w[199][166] = 5'b01111; w[199][167] = 5'b01111; w[199][168] = 5'b01111; w[199][169] = 5'b01111; w[199][170] = 5'b01111; w[199][171] = 5'b01111; w[199][172] = 5'b00000; w[199][173] = 5'b00000; w[199][174] = 5'b10000; w[199][175] = 5'b10000; w[199][176] = 5'b10000; w[199][177] = 5'b00000; w[199][178] = 5'b01111; w[199][179] = 5'b01111; w[199][180] = 5'b01111; w[199][181] = 5'b01111; w[199][182] = 5'b01111; w[199][183] = 5'b01111; w[199][184] = 5'b01111; w[199][185] = 5'b01111; w[199][186] = 5'b01111; w[199][187] = 5'b01111; w[199][188] = 5'b01111; w[199][189] = 5'b01111; w[199][190] = 5'b01111; w[199][191] = 5'b01111; w[199][192] = 5'b01111; w[199][193] = 5'b01111; w[199][194] = 5'b01111; w[199][195] = 5'b01111; w[199][196] = 5'b01111; w[199][197] = 5'b01111; w[199][198] = 5'b01111; w[199][199] = 5'b00000; w[199][200] = 5'b01111; w[199][201] = 5'b01111; w[199][202] = 5'b01111; w[199][203] = 5'b01111; w[199][204] = 5'b01111; w[199][205] = 5'b01111; w[199][206] = 5'b01111; w[199][207] = 5'b01111; w[199][208] = 5'b01111; w[199][209] = 5'b01111; 
w[200][0] = 5'b01111; w[200][1] = 5'b01111; w[200][2] = 5'b01111; w[200][3] = 5'b01111; w[200][4] = 5'b01111; w[200][5] = 5'b01111; w[200][6] = 5'b01111; w[200][7] = 5'b01111; w[200][8] = 5'b01111; w[200][9] = 5'b01111; w[200][10] = 5'b01111; w[200][11] = 5'b01111; w[200][12] = 5'b01111; w[200][13] = 5'b01111; w[200][14] = 5'b01111; w[200][15] = 5'b01111; w[200][16] = 5'b01111; w[200][17] = 5'b01111; w[200][18] = 5'b01111; w[200][19] = 5'b01111; w[200][20] = 5'b01111; w[200][21] = 5'b01111; w[200][22] = 5'b01111; w[200][23] = 5'b01111; w[200][24] = 5'b01111; w[200][25] = 5'b01111; w[200][26] = 5'b01111; w[200][27] = 5'b01111; w[200][28] = 5'b01111; w[200][29] = 5'b01111; w[200][30] = 5'b01111; w[200][31] = 5'b00000; w[200][32] = 5'b10000; w[200][33] = 5'b10000; w[200][34] = 5'b10000; w[200][35] = 5'b10000; w[200][36] = 5'b10000; w[200][37] = 5'b10000; w[200][38] = 5'b00000; w[200][39] = 5'b01111; w[200][40] = 5'b01111; w[200][41] = 5'b01111; w[200][42] = 5'b01111; w[200][43] = 5'b01111; w[200][44] = 5'b01111; w[200][45] = 5'b10000; w[200][46] = 5'b10000; w[200][47] = 5'b10000; w[200][48] = 5'b10000; w[200][49] = 5'b10000; w[200][50] = 5'b10000; w[200][51] = 5'b10000; w[200][52] = 5'b10000; w[200][53] = 5'b01111; w[200][54] = 5'b01111; w[200][55] = 5'b01111; w[200][56] = 5'b01111; w[200][57] = 5'b01111; w[200][58] = 5'b01111; w[200][59] = 5'b00000; w[200][60] = 5'b00000; w[200][61] = 5'b01111; w[200][62] = 5'b10000; w[200][63] = 5'b00000; w[200][64] = 5'b01111; w[200][65] = 5'b00000; w[200][66] = 5'b00000; w[200][67] = 5'b01111; w[200][68] = 5'b01111; w[200][69] = 5'b01111; w[200][70] = 5'b01111; w[200][71] = 5'b01111; w[200][72] = 5'b01111; w[200][73] = 5'b00000; w[200][74] = 5'b01111; w[200][75] = 5'b01111; w[200][76] = 5'b10000; w[200][77] = 5'b00000; w[200][78] = 5'b01111; w[200][79] = 5'b01111; w[200][80] = 5'b00000; w[200][81] = 5'b01111; w[200][82] = 5'b01111; w[200][83] = 5'b01111; w[200][84] = 5'b01111; w[200][85] = 5'b01111; w[200][86] = 5'b01111; w[200][87] = 5'b00000; w[200][88] = 5'b01111; w[200][89] = 5'b01111; w[200][90] = 5'b10000; w[200][91] = 5'b10000; w[200][92] = 5'b01111; w[200][93] = 5'b01111; w[200][94] = 5'b01111; w[200][95] = 5'b01111; w[200][96] = 5'b01111; w[200][97] = 5'b01111; w[200][98] = 5'b01111; w[200][99] = 5'b01111; w[200][100] = 5'b01111; w[200][101] = 5'b00000; w[200][102] = 5'b01111; w[200][103] = 5'b01111; w[200][104] = 5'b10000; w[200][105] = 5'b10000; w[200][106] = 5'b01111; w[200][107] = 5'b00000; w[200][108] = 5'b00000; w[200][109] = 5'b01111; w[200][110] = 5'b01111; w[200][111] = 5'b01111; w[200][112] = 5'b01111; w[200][113] = 5'b01111; w[200][114] = 5'b01111; w[200][115] = 5'b00000; w[200][116] = 5'b01111; w[200][117] = 5'b01111; w[200][118] = 5'b10000; w[200][119] = 5'b10000; w[200][120] = 5'b00000; w[200][121] = 5'b00000; w[200][122] = 5'b00000; w[200][123] = 5'b01111; w[200][124] = 5'b01111; w[200][125] = 5'b01111; w[200][126] = 5'b01111; w[200][127] = 5'b01111; w[200][128] = 5'b01111; w[200][129] = 5'b00000; w[200][130] = 5'b01111; w[200][131] = 5'b01111; w[200][132] = 5'b00000; w[200][133] = 5'b10000; w[200][134] = 5'b01111; w[200][135] = 5'b01111; w[200][136] = 5'b00000; w[200][137] = 5'b01111; w[200][138] = 5'b01111; w[200][139] = 5'b01111; w[200][140] = 5'b01111; w[200][141] = 5'b01111; w[200][142] = 5'b01111; w[200][143] = 5'b00000; w[200][144] = 5'b00000; w[200][145] = 5'b01111; w[200][146] = 5'b00000; w[200][147] = 5'b10000; w[200][148] = 5'b01111; w[200][149] = 5'b00000; w[200][150] = 5'b00000; w[200][151] = 5'b01111; w[200][152] = 5'b01111; w[200][153] = 5'b01111; w[200][154] = 5'b01111; w[200][155] = 5'b01111; w[200][156] = 5'b01111; w[200][157] = 5'b00000; w[200][158] = 5'b00000; w[200][159] = 5'b00000; w[200][160] = 5'b10000; w[200][161] = 5'b10000; w[200][162] = 5'b10000; w[200][163] = 5'b00000; w[200][164] = 5'b00000; w[200][165] = 5'b01111; w[200][166] = 5'b01111; w[200][167] = 5'b01111; w[200][168] = 5'b01111; w[200][169] = 5'b01111; w[200][170] = 5'b01111; w[200][171] = 5'b01111; w[200][172] = 5'b00000; w[200][173] = 5'b00000; w[200][174] = 5'b10000; w[200][175] = 5'b10000; w[200][176] = 5'b10000; w[200][177] = 5'b00000; w[200][178] = 5'b01111; w[200][179] = 5'b01111; w[200][180] = 5'b01111; w[200][181] = 5'b01111; w[200][182] = 5'b01111; w[200][183] = 5'b01111; w[200][184] = 5'b01111; w[200][185] = 5'b01111; w[200][186] = 5'b01111; w[200][187] = 5'b01111; w[200][188] = 5'b01111; w[200][189] = 5'b01111; w[200][190] = 5'b01111; w[200][191] = 5'b01111; w[200][192] = 5'b01111; w[200][193] = 5'b01111; w[200][194] = 5'b01111; w[200][195] = 5'b01111; w[200][196] = 5'b01111; w[200][197] = 5'b01111; w[200][198] = 5'b01111; w[200][199] = 5'b01111; w[200][200] = 5'b00000; w[200][201] = 5'b01111; w[200][202] = 5'b01111; w[200][203] = 5'b01111; w[200][204] = 5'b01111; w[200][205] = 5'b01111; w[200][206] = 5'b01111; w[200][207] = 5'b01111; w[200][208] = 5'b01111; w[200][209] = 5'b01111; 
w[201][0] = 5'b01111; w[201][1] = 5'b01111; w[201][2] = 5'b01111; w[201][3] = 5'b01111; w[201][4] = 5'b01111; w[201][5] = 5'b01111; w[201][6] = 5'b01111; w[201][7] = 5'b01111; w[201][8] = 5'b01111; w[201][9] = 5'b01111; w[201][10] = 5'b01111; w[201][11] = 5'b01111; w[201][12] = 5'b01111; w[201][13] = 5'b01111; w[201][14] = 5'b01111; w[201][15] = 5'b01111; w[201][16] = 5'b01111; w[201][17] = 5'b01111; w[201][18] = 5'b01111; w[201][19] = 5'b01111; w[201][20] = 5'b01111; w[201][21] = 5'b01111; w[201][22] = 5'b01111; w[201][23] = 5'b01111; w[201][24] = 5'b01111; w[201][25] = 5'b01111; w[201][26] = 5'b01111; w[201][27] = 5'b01111; w[201][28] = 5'b01111; w[201][29] = 5'b01111; w[201][30] = 5'b01111; w[201][31] = 5'b00000; w[201][32] = 5'b10000; w[201][33] = 5'b10000; w[201][34] = 5'b10000; w[201][35] = 5'b10000; w[201][36] = 5'b10000; w[201][37] = 5'b10000; w[201][38] = 5'b00000; w[201][39] = 5'b01111; w[201][40] = 5'b01111; w[201][41] = 5'b01111; w[201][42] = 5'b01111; w[201][43] = 5'b01111; w[201][44] = 5'b01111; w[201][45] = 5'b10000; w[201][46] = 5'b10000; w[201][47] = 5'b10000; w[201][48] = 5'b10000; w[201][49] = 5'b10000; w[201][50] = 5'b10000; w[201][51] = 5'b10000; w[201][52] = 5'b10000; w[201][53] = 5'b01111; w[201][54] = 5'b01111; w[201][55] = 5'b01111; w[201][56] = 5'b01111; w[201][57] = 5'b01111; w[201][58] = 5'b01111; w[201][59] = 5'b00000; w[201][60] = 5'b00000; w[201][61] = 5'b01111; w[201][62] = 5'b10000; w[201][63] = 5'b00000; w[201][64] = 5'b01111; w[201][65] = 5'b00000; w[201][66] = 5'b00000; w[201][67] = 5'b01111; w[201][68] = 5'b01111; w[201][69] = 5'b01111; w[201][70] = 5'b01111; w[201][71] = 5'b01111; w[201][72] = 5'b01111; w[201][73] = 5'b00000; w[201][74] = 5'b01111; w[201][75] = 5'b01111; w[201][76] = 5'b10000; w[201][77] = 5'b00000; w[201][78] = 5'b01111; w[201][79] = 5'b01111; w[201][80] = 5'b00000; w[201][81] = 5'b01111; w[201][82] = 5'b01111; w[201][83] = 5'b01111; w[201][84] = 5'b01111; w[201][85] = 5'b01111; w[201][86] = 5'b01111; w[201][87] = 5'b00000; w[201][88] = 5'b01111; w[201][89] = 5'b01111; w[201][90] = 5'b10000; w[201][91] = 5'b10000; w[201][92] = 5'b01111; w[201][93] = 5'b01111; w[201][94] = 5'b01111; w[201][95] = 5'b01111; w[201][96] = 5'b01111; w[201][97] = 5'b01111; w[201][98] = 5'b01111; w[201][99] = 5'b01111; w[201][100] = 5'b01111; w[201][101] = 5'b00000; w[201][102] = 5'b01111; w[201][103] = 5'b01111; w[201][104] = 5'b10000; w[201][105] = 5'b10000; w[201][106] = 5'b01111; w[201][107] = 5'b00000; w[201][108] = 5'b00000; w[201][109] = 5'b01111; w[201][110] = 5'b01111; w[201][111] = 5'b01111; w[201][112] = 5'b01111; w[201][113] = 5'b01111; w[201][114] = 5'b01111; w[201][115] = 5'b00000; w[201][116] = 5'b01111; w[201][117] = 5'b01111; w[201][118] = 5'b10000; w[201][119] = 5'b10000; w[201][120] = 5'b00000; w[201][121] = 5'b00000; w[201][122] = 5'b00000; w[201][123] = 5'b01111; w[201][124] = 5'b01111; w[201][125] = 5'b01111; w[201][126] = 5'b01111; w[201][127] = 5'b01111; w[201][128] = 5'b01111; w[201][129] = 5'b00000; w[201][130] = 5'b01111; w[201][131] = 5'b01111; w[201][132] = 5'b00000; w[201][133] = 5'b10000; w[201][134] = 5'b01111; w[201][135] = 5'b01111; w[201][136] = 5'b00000; w[201][137] = 5'b01111; w[201][138] = 5'b01111; w[201][139] = 5'b01111; w[201][140] = 5'b01111; w[201][141] = 5'b01111; w[201][142] = 5'b01111; w[201][143] = 5'b00000; w[201][144] = 5'b00000; w[201][145] = 5'b01111; w[201][146] = 5'b00000; w[201][147] = 5'b10000; w[201][148] = 5'b01111; w[201][149] = 5'b00000; w[201][150] = 5'b00000; w[201][151] = 5'b01111; w[201][152] = 5'b01111; w[201][153] = 5'b01111; w[201][154] = 5'b01111; w[201][155] = 5'b01111; w[201][156] = 5'b01111; w[201][157] = 5'b00000; w[201][158] = 5'b00000; w[201][159] = 5'b00000; w[201][160] = 5'b10000; w[201][161] = 5'b10000; w[201][162] = 5'b10000; w[201][163] = 5'b00000; w[201][164] = 5'b00000; w[201][165] = 5'b01111; w[201][166] = 5'b01111; w[201][167] = 5'b01111; w[201][168] = 5'b01111; w[201][169] = 5'b01111; w[201][170] = 5'b01111; w[201][171] = 5'b01111; w[201][172] = 5'b00000; w[201][173] = 5'b00000; w[201][174] = 5'b10000; w[201][175] = 5'b10000; w[201][176] = 5'b10000; w[201][177] = 5'b00000; w[201][178] = 5'b01111; w[201][179] = 5'b01111; w[201][180] = 5'b01111; w[201][181] = 5'b01111; w[201][182] = 5'b01111; w[201][183] = 5'b01111; w[201][184] = 5'b01111; w[201][185] = 5'b01111; w[201][186] = 5'b01111; w[201][187] = 5'b01111; w[201][188] = 5'b01111; w[201][189] = 5'b01111; w[201][190] = 5'b01111; w[201][191] = 5'b01111; w[201][192] = 5'b01111; w[201][193] = 5'b01111; w[201][194] = 5'b01111; w[201][195] = 5'b01111; w[201][196] = 5'b01111; w[201][197] = 5'b01111; w[201][198] = 5'b01111; w[201][199] = 5'b01111; w[201][200] = 5'b01111; w[201][201] = 5'b00000; w[201][202] = 5'b01111; w[201][203] = 5'b01111; w[201][204] = 5'b01111; w[201][205] = 5'b01111; w[201][206] = 5'b01111; w[201][207] = 5'b01111; w[201][208] = 5'b01111; w[201][209] = 5'b01111; 
w[202][0] = 5'b01111; w[202][1] = 5'b01111; w[202][2] = 5'b01111; w[202][3] = 5'b01111; w[202][4] = 5'b01111; w[202][5] = 5'b01111; w[202][6] = 5'b01111; w[202][7] = 5'b01111; w[202][8] = 5'b01111; w[202][9] = 5'b01111; w[202][10] = 5'b01111; w[202][11] = 5'b01111; w[202][12] = 5'b01111; w[202][13] = 5'b01111; w[202][14] = 5'b01111; w[202][15] = 5'b01111; w[202][16] = 5'b01111; w[202][17] = 5'b01111; w[202][18] = 5'b01111; w[202][19] = 5'b01111; w[202][20] = 5'b01111; w[202][21] = 5'b01111; w[202][22] = 5'b01111; w[202][23] = 5'b01111; w[202][24] = 5'b01111; w[202][25] = 5'b01111; w[202][26] = 5'b01111; w[202][27] = 5'b01111; w[202][28] = 5'b01111; w[202][29] = 5'b01111; w[202][30] = 5'b01111; w[202][31] = 5'b00000; w[202][32] = 5'b10000; w[202][33] = 5'b10000; w[202][34] = 5'b10000; w[202][35] = 5'b10000; w[202][36] = 5'b10000; w[202][37] = 5'b10000; w[202][38] = 5'b00000; w[202][39] = 5'b01111; w[202][40] = 5'b01111; w[202][41] = 5'b01111; w[202][42] = 5'b01111; w[202][43] = 5'b01111; w[202][44] = 5'b01111; w[202][45] = 5'b10000; w[202][46] = 5'b10000; w[202][47] = 5'b10000; w[202][48] = 5'b10000; w[202][49] = 5'b10000; w[202][50] = 5'b10000; w[202][51] = 5'b10000; w[202][52] = 5'b10000; w[202][53] = 5'b01111; w[202][54] = 5'b01111; w[202][55] = 5'b01111; w[202][56] = 5'b01111; w[202][57] = 5'b01111; w[202][58] = 5'b01111; w[202][59] = 5'b00000; w[202][60] = 5'b00000; w[202][61] = 5'b01111; w[202][62] = 5'b10000; w[202][63] = 5'b00000; w[202][64] = 5'b01111; w[202][65] = 5'b00000; w[202][66] = 5'b00000; w[202][67] = 5'b01111; w[202][68] = 5'b01111; w[202][69] = 5'b01111; w[202][70] = 5'b01111; w[202][71] = 5'b01111; w[202][72] = 5'b01111; w[202][73] = 5'b00000; w[202][74] = 5'b01111; w[202][75] = 5'b01111; w[202][76] = 5'b10000; w[202][77] = 5'b00000; w[202][78] = 5'b01111; w[202][79] = 5'b01111; w[202][80] = 5'b00000; w[202][81] = 5'b01111; w[202][82] = 5'b01111; w[202][83] = 5'b01111; w[202][84] = 5'b01111; w[202][85] = 5'b01111; w[202][86] = 5'b01111; w[202][87] = 5'b00000; w[202][88] = 5'b01111; w[202][89] = 5'b01111; w[202][90] = 5'b10000; w[202][91] = 5'b10000; w[202][92] = 5'b01111; w[202][93] = 5'b01111; w[202][94] = 5'b01111; w[202][95] = 5'b01111; w[202][96] = 5'b01111; w[202][97] = 5'b01111; w[202][98] = 5'b01111; w[202][99] = 5'b01111; w[202][100] = 5'b01111; w[202][101] = 5'b00000; w[202][102] = 5'b01111; w[202][103] = 5'b01111; w[202][104] = 5'b10000; w[202][105] = 5'b10000; w[202][106] = 5'b01111; w[202][107] = 5'b00000; w[202][108] = 5'b00000; w[202][109] = 5'b01111; w[202][110] = 5'b01111; w[202][111] = 5'b01111; w[202][112] = 5'b01111; w[202][113] = 5'b01111; w[202][114] = 5'b01111; w[202][115] = 5'b00000; w[202][116] = 5'b01111; w[202][117] = 5'b01111; w[202][118] = 5'b10000; w[202][119] = 5'b10000; w[202][120] = 5'b00000; w[202][121] = 5'b00000; w[202][122] = 5'b00000; w[202][123] = 5'b01111; w[202][124] = 5'b01111; w[202][125] = 5'b01111; w[202][126] = 5'b01111; w[202][127] = 5'b01111; w[202][128] = 5'b01111; w[202][129] = 5'b00000; w[202][130] = 5'b01111; w[202][131] = 5'b01111; w[202][132] = 5'b00000; w[202][133] = 5'b10000; w[202][134] = 5'b01111; w[202][135] = 5'b01111; w[202][136] = 5'b00000; w[202][137] = 5'b01111; w[202][138] = 5'b01111; w[202][139] = 5'b01111; w[202][140] = 5'b01111; w[202][141] = 5'b01111; w[202][142] = 5'b01111; w[202][143] = 5'b00000; w[202][144] = 5'b00000; w[202][145] = 5'b01111; w[202][146] = 5'b00000; w[202][147] = 5'b10000; w[202][148] = 5'b01111; w[202][149] = 5'b00000; w[202][150] = 5'b00000; w[202][151] = 5'b01111; w[202][152] = 5'b01111; w[202][153] = 5'b01111; w[202][154] = 5'b01111; w[202][155] = 5'b01111; w[202][156] = 5'b01111; w[202][157] = 5'b00000; w[202][158] = 5'b00000; w[202][159] = 5'b00000; w[202][160] = 5'b10000; w[202][161] = 5'b10000; w[202][162] = 5'b10000; w[202][163] = 5'b00000; w[202][164] = 5'b00000; w[202][165] = 5'b01111; w[202][166] = 5'b01111; w[202][167] = 5'b01111; w[202][168] = 5'b01111; w[202][169] = 5'b01111; w[202][170] = 5'b01111; w[202][171] = 5'b01111; w[202][172] = 5'b00000; w[202][173] = 5'b00000; w[202][174] = 5'b10000; w[202][175] = 5'b10000; w[202][176] = 5'b10000; w[202][177] = 5'b00000; w[202][178] = 5'b01111; w[202][179] = 5'b01111; w[202][180] = 5'b01111; w[202][181] = 5'b01111; w[202][182] = 5'b01111; w[202][183] = 5'b01111; w[202][184] = 5'b01111; w[202][185] = 5'b01111; w[202][186] = 5'b01111; w[202][187] = 5'b01111; w[202][188] = 5'b01111; w[202][189] = 5'b01111; w[202][190] = 5'b01111; w[202][191] = 5'b01111; w[202][192] = 5'b01111; w[202][193] = 5'b01111; w[202][194] = 5'b01111; w[202][195] = 5'b01111; w[202][196] = 5'b01111; w[202][197] = 5'b01111; w[202][198] = 5'b01111; w[202][199] = 5'b01111; w[202][200] = 5'b01111; w[202][201] = 5'b01111; w[202][202] = 5'b00000; w[202][203] = 5'b01111; w[202][204] = 5'b01111; w[202][205] = 5'b01111; w[202][206] = 5'b01111; w[202][207] = 5'b01111; w[202][208] = 5'b01111; w[202][209] = 5'b01111; 
w[203][0] = 5'b01111; w[203][1] = 5'b01111; w[203][2] = 5'b01111; w[203][3] = 5'b01111; w[203][4] = 5'b01111; w[203][5] = 5'b01111; w[203][6] = 5'b01111; w[203][7] = 5'b01111; w[203][8] = 5'b01111; w[203][9] = 5'b01111; w[203][10] = 5'b01111; w[203][11] = 5'b01111; w[203][12] = 5'b01111; w[203][13] = 5'b01111; w[203][14] = 5'b01111; w[203][15] = 5'b01111; w[203][16] = 5'b01111; w[203][17] = 5'b01111; w[203][18] = 5'b01111; w[203][19] = 5'b01111; w[203][20] = 5'b01111; w[203][21] = 5'b01111; w[203][22] = 5'b01111; w[203][23] = 5'b01111; w[203][24] = 5'b01111; w[203][25] = 5'b01111; w[203][26] = 5'b01111; w[203][27] = 5'b01111; w[203][28] = 5'b01111; w[203][29] = 5'b01111; w[203][30] = 5'b01111; w[203][31] = 5'b00000; w[203][32] = 5'b10000; w[203][33] = 5'b10000; w[203][34] = 5'b10000; w[203][35] = 5'b10000; w[203][36] = 5'b10000; w[203][37] = 5'b10000; w[203][38] = 5'b00000; w[203][39] = 5'b01111; w[203][40] = 5'b01111; w[203][41] = 5'b01111; w[203][42] = 5'b01111; w[203][43] = 5'b01111; w[203][44] = 5'b01111; w[203][45] = 5'b10000; w[203][46] = 5'b10000; w[203][47] = 5'b10000; w[203][48] = 5'b10000; w[203][49] = 5'b10000; w[203][50] = 5'b10000; w[203][51] = 5'b10000; w[203][52] = 5'b10000; w[203][53] = 5'b01111; w[203][54] = 5'b01111; w[203][55] = 5'b01111; w[203][56] = 5'b01111; w[203][57] = 5'b01111; w[203][58] = 5'b01111; w[203][59] = 5'b00000; w[203][60] = 5'b00000; w[203][61] = 5'b01111; w[203][62] = 5'b10000; w[203][63] = 5'b00000; w[203][64] = 5'b01111; w[203][65] = 5'b00000; w[203][66] = 5'b00000; w[203][67] = 5'b01111; w[203][68] = 5'b01111; w[203][69] = 5'b01111; w[203][70] = 5'b01111; w[203][71] = 5'b01111; w[203][72] = 5'b01111; w[203][73] = 5'b00000; w[203][74] = 5'b01111; w[203][75] = 5'b01111; w[203][76] = 5'b10000; w[203][77] = 5'b00000; w[203][78] = 5'b01111; w[203][79] = 5'b01111; w[203][80] = 5'b00000; w[203][81] = 5'b01111; w[203][82] = 5'b01111; w[203][83] = 5'b01111; w[203][84] = 5'b01111; w[203][85] = 5'b01111; w[203][86] = 5'b01111; w[203][87] = 5'b00000; w[203][88] = 5'b01111; w[203][89] = 5'b01111; w[203][90] = 5'b10000; w[203][91] = 5'b10000; w[203][92] = 5'b01111; w[203][93] = 5'b01111; w[203][94] = 5'b01111; w[203][95] = 5'b01111; w[203][96] = 5'b01111; w[203][97] = 5'b01111; w[203][98] = 5'b01111; w[203][99] = 5'b01111; w[203][100] = 5'b01111; w[203][101] = 5'b00000; w[203][102] = 5'b01111; w[203][103] = 5'b01111; w[203][104] = 5'b10000; w[203][105] = 5'b10000; w[203][106] = 5'b01111; w[203][107] = 5'b00000; w[203][108] = 5'b00000; w[203][109] = 5'b01111; w[203][110] = 5'b01111; w[203][111] = 5'b01111; w[203][112] = 5'b01111; w[203][113] = 5'b01111; w[203][114] = 5'b01111; w[203][115] = 5'b00000; w[203][116] = 5'b01111; w[203][117] = 5'b01111; w[203][118] = 5'b10000; w[203][119] = 5'b10000; w[203][120] = 5'b00000; w[203][121] = 5'b00000; w[203][122] = 5'b00000; w[203][123] = 5'b01111; w[203][124] = 5'b01111; w[203][125] = 5'b01111; w[203][126] = 5'b01111; w[203][127] = 5'b01111; w[203][128] = 5'b01111; w[203][129] = 5'b00000; w[203][130] = 5'b01111; w[203][131] = 5'b01111; w[203][132] = 5'b00000; w[203][133] = 5'b10000; w[203][134] = 5'b01111; w[203][135] = 5'b01111; w[203][136] = 5'b00000; w[203][137] = 5'b01111; w[203][138] = 5'b01111; w[203][139] = 5'b01111; w[203][140] = 5'b01111; w[203][141] = 5'b01111; w[203][142] = 5'b01111; w[203][143] = 5'b00000; w[203][144] = 5'b00000; w[203][145] = 5'b01111; w[203][146] = 5'b00000; w[203][147] = 5'b10000; w[203][148] = 5'b01111; w[203][149] = 5'b00000; w[203][150] = 5'b00000; w[203][151] = 5'b01111; w[203][152] = 5'b01111; w[203][153] = 5'b01111; w[203][154] = 5'b01111; w[203][155] = 5'b01111; w[203][156] = 5'b01111; w[203][157] = 5'b00000; w[203][158] = 5'b00000; w[203][159] = 5'b00000; w[203][160] = 5'b10000; w[203][161] = 5'b10000; w[203][162] = 5'b10000; w[203][163] = 5'b00000; w[203][164] = 5'b00000; w[203][165] = 5'b01111; w[203][166] = 5'b01111; w[203][167] = 5'b01111; w[203][168] = 5'b01111; w[203][169] = 5'b01111; w[203][170] = 5'b01111; w[203][171] = 5'b01111; w[203][172] = 5'b00000; w[203][173] = 5'b00000; w[203][174] = 5'b10000; w[203][175] = 5'b10000; w[203][176] = 5'b10000; w[203][177] = 5'b00000; w[203][178] = 5'b01111; w[203][179] = 5'b01111; w[203][180] = 5'b01111; w[203][181] = 5'b01111; w[203][182] = 5'b01111; w[203][183] = 5'b01111; w[203][184] = 5'b01111; w[203][185] = 5'b01111; w[203][186] = 5'b01111; w[203][187] = 5'b01111; w[203][188] = 5'b01111; w[203][189] = 5'b01111; w[203][190] = 5'b01111; w[203][191] = 5'b01111; w[203][192] = 5'b01111; w[203][193] = 5'b01111; w[203][194] = 5'b01111; w[203][195] = 5'b01111; w[203][196] = 5'b01111; w[203][197] = 5'b01111; w[203][198] = 5'b01111; w[203][199] = 5'b01111; w[203][200] = 5'b01111; w[203][201] = 5'b01111; w[203][202] = 5'b01111; w[203][203] = 5'b00000; w[203][204] = 5'b01111; w[203][205] = 5'b01111; w[203][206] = 5'b01111; w[203][207] = 5'b01111; w[203][208] = 5'b01111; w[203][209] = 5'b01111; 
w[204][0] = 5'b01111; w[204][1] = 5'b01111; w[204][2] = 5'b01111; w[204][3] = 5'b01111; w[204][4] = 5'b01111; w[204][5] = 5'b01111; w[204][6] = 5'b01111; w[204][7] = 5'b01111; w[204][8] = 5'b01111; w[204][9] = 5'b01111; w[204][10] = 5'b01111; w[204][11] = 5'b01111; w[204][12] = 5'b01111; w[204][13] = 5'b01111; w[204][14] = 5'b01111; w[204][15] = 5'b01111; w[204][16] = 5'b01111; w[204][17] = 5'b01111; w[204][18] = 5'b01111; w[204][19] = 5'b01111; w[204][20] = 5'b01111; w[204][21] = 5'b01111; w[204][22] = 5'b01111; w[204][23] = 5'b01111; w[204][24] = 5'b01111; w[204][25] = 5'b01111; w[204][26] = 5'b01111; w[204][27] = 5'b01111; w[204][28] = 5'b01111; w[204][29] = 5'b01111; w[204][30] = 5'b01111; w[204][31] = 5'b00000; w[204][32] = 5'b10000; w[204][33] = 5'b10000; w[204][34] = 5'b10000; w[204][35] = 5'b10000; w[204][36] = 5'b10000; w[204][37] = 5'b10000; w[204][38] = 5'b00000; w[204][39] = 5'b01111; w[204][40] = 5'b01111; w[204][41] = 5'b01111; w[204][42] = 5'b01111; w[204][43] = 5'b01111; w[204][44] = 5'b01111; w[204][45] = 5'b10000; w[204][46] = 5'b10000; w[204][47] = 5'b10000; w[204][48] = 5'b10000; w[204][49] = 5'b10000; w[204][50] = 5'b10000; w[204][51] = 5'b10000; w[204][52] = 5'b10000; w[204][53] = 5'b01111; w[204][54] = 5'b01111; w[204][55] = 5'b01111; w[204][56] = 5'b01111; w[204][57] = 5'b01111; w[204][58] = 5'b01111; w[204][59] = 5'b00000; w[204][60] = 5'b00000; w[204][61] = 5'b01111; w[204][62] = 5'b10000; w[204][63] = 5'b00000; w[204][64] = 5'b01111; w[204][65] = 5'b00000; w[204][66] = 5'b00000; w[204][67] = 5'b01111; w[204][68] = 5'b01111; w[204][69] = 5'b01111; w[204][70] = 5'b01111; w[204][71] = 5'b01111; w[204][72] = 5'b01111; w[204][73] = 5'b00000; w[204][74] = 5'b01111; w[204][75] = 5'b01111; w[204][76] = 5'b10000; w[204][77] = 5'b00000; w[204][78] = 5'b01111; w[204][79] = 5'b01111; w[204][80] = 5'b00000; w[204][81] = 5'b01111; w[204][82] = 5'b01111; w[204][83] = 5'b01111; w[204][84] = 5'b01111; w[204][85] = 5'b01111; w[204][86] = 5'b01111; w[204][87] = 5'b00000; w[204][88] = 5'b01111; w[204][89] = 5'b01111; w[204][90] = 5'b10000; w[204][91] = 5'b10000; w[204][92] = 5'b01111; w[204][93] = 5'b01111; w[204][94] = 5'b01111; w[204][95] = 5'b01111; w[204][96] = 5'b01111; w[204][97] = 5'b01111; w[204][98] = 5'b01111; w[204][99] = 5'b01111; w[204][100] = 5'b01111; w[204][101] = 5'b00000; w[204][102] = 5'b01111; w[204][103] = 5'b01111; w[204][104] = 5'b10000; w[204][105] = 5'b10000; w[204][106] = 5'b01111; w[204][107] = 5'b00000; w[204][108] = 5'b00000; w[204][109] = 5'b01111; w[204][110] = 5'b01111; w[204][111] = 5'b01111; w[204][112] = 5'b01111; w[204][113] = 5'b01111; w[204][114] = 5'b01111; w[204][115] = 5'b00000; w[204][116] = 5'b01111; w[204][117] = 5'b01111; w[204][118] = 5'b10000; w[204][119] = 5'b10000; w[204][120] = 5'b00000; w[204][121] = 5'b00000; w[204][122] = 5'b00000; w[204][123] = 5'b01111; w[204][124] = 5'b01111; w[204][125] = 5'b01111; w[204][126] = 5'b01111; w[204][127] = 5'b01111; w[204][128] = 5'b01111; w[204][129] = 5'b00000; w[204][130] = 5'b01111; w[204][131] = 5'b01111; w[204][132] = 5'b00000; w[204][133] = 5'b10000; w[204][134] = 5'b01111; w[204][135] = 5'b01111; w[204][136] = 5'b00000; w[204][137] = 5'b01111; w[204][138] = 5'b01111; w[204][139] = 5'b01111; w[204][140] = 5'b01111; w[204][141] = 5'b01111; w[204][142] = 5'b01111; w[204][143] = 5'b00000; w[204][144] = 5'b00000; w[204][145] = 5'b01111; w[204][146] = 5'b00000; w[204][147] = 5'b10000; w[204][148] = 5'b01111; w[204][149] = 5'b00000; w[204][150] = 5'b00000; w[204][151] = 5'b01111; w[204][152] = 5'b01111; w[204][153] = 5'b01111; w[204][154] = 5'b01111; w[204][155] = 5'b01111; w[204][156] = 5'b01111; w[204][157] = 5'b00000; w[204][158] = 5'b00000; w[204][159] = 5'b00000; w[204][160] = 5'b10000; w[204][161] = 5'b10000; w[204][162] = 5'b10000; w[204][163] = 5'b00000; w[204][164] = 5'b00000; w[204][165] = 5'b01111; w[204][166] = 5'b01111; w[204][167] = 5'b01111; w[204][168] = 5'b01111; w[204][169] = 5'b01111; w[204][170] = 5'b01111; w[204][171] = 5'b01111; w[204][172] = 5'b00000; w[204][173] = 5'b00000; w[204][174] = 5'b10000; w[204][175] = 5'b10000; w[204][176] = 5'b10000; w[204][177] = 5'b00000; w[204][178] = 5'b01111; w[204][179] = 5'b01111; w[204][180] = 5'b01111; w[204][181] = 5'b01111; w[204][182] = 5'b01111; w[204][183] = 5'b01111; w[204][184] = 5'b01111; w[204][185] = 5'b01111; w[204][186] = 5'b01111; w[204][187] = 5'b01111; w[204][188] = 5'b01111; w[204][189] = 5'b01111; w[204][190] = 5'b01111; w[204][191] = 5'b01111; w[204][192] = 5'b01111; w[204][193] = 5'b01111; w[204][194] = 5'b01111; w[204][195] = 5'b01111; w[204][196] = 5'b01111; w[204][197] = 5'b01111; w[204][198] = 5'b01111; w[204][199] = 5'b01111; w[204][200] = 5'b01111; w[204][201] = 5'b01111; w[204][202] = 5'b01111; w[204][203] = 5'b01111; w[204][204] = 5'b00000; w[204][205] = 5'b01111; w[204][206] = 5'b01111; w[204][207] = 5'b01111; w[204][208] = 5'b01111; w[204][209] = 5'b01111; 
w[205][0] = 5'b01111; w[205][1] = 5'b01111; w[205][2] = 5'b01111; w[205][3] = 5'b01111; w[205][4] = 5'b01111; w[205][5] = 5'b01111; w[205][6] = 5'b01111; w[205][7] = 5'b01111; w[205][8] = 5'b01111; w[205][9] = 5'b01111; w[205][10] = 5'b01111; w[205][11] = 5'b01111; w[205][12] = 5'b01111; w[205][13] = 5'b01111; w[205][14] = 5'b01111; w[205][15] = 5'b01111; w[205][16] = 5'b01111; w[205][17] = 5'b01111; w[205][18] = 5'b01111; w[205][19] = 5'b01111; w[205][20] = 5'b01111; w[205][21] = 5'b01111; w[205][22] = 5'b01111; w[205][23] = 5'b01111; w[205][24] = 5'b01111; w[205][25] = 5'b01111; w[205][26] = 5'b01111; w[205][27] = 5'b01111; w[205][28] = 5'b01111; w[205][29] = 5'b01111; w[205][30] = 5'b01111; w[205][31] = 5'b00000; w[205][32] = 5'b10000; w[205][33] = 5'b10000; w[205][34] = 5'b10000; w[205][35] = 5'b10000; w[205][36] = 5'b10000; w[205][37] = 5'b10000; w[205][38] = 5'b00000; w[205][39] = 5'b01111; w[205][40] = 5'b01111; w[205][41] = 5'b01111; w[205][42] = 5'b01111; w[205][43] = 5'b01111; w[205][44] = 5'b01111; w[205][45] = 5'b10000; w[205][46] = 5'b10000; w[205][47] = 5'b10000; w[205][48] = 5'b10000; w[205][49] = 5'b10000; w[205][50] = 5'b10000; w[205][51] = 5'b10000; w[205][52] = 5'b10000; w[205][53] = 5'b01111; w[205][54] = 5'b01111; w[205][55] = 5'b01111; w[205][56] = 5'b01111; w[205][57] = 5'b01111; w[205][58] = 5'b01111; w[205][59] = 5'b00000; w[205][60] = 5'b00000; w[205][61] = 5'b01111; w[205][62] = 5'b10000; w[205][63] = 5'b00000; w[205][64] = 5'b01111; w[205][65] = 5'b00000; w[205][66] = 5'b00000; w[205][67] = 5'b01111; w[205][68] = 5'b01111; w[205][69] = 5'b01111; w[205][70] = 5'b01111; w[205][71] = 5'b01111; w[205][72] = 5'b01111; w[205][73] = 5'b00000; w[205][74] = 5'b01111; w[205][75] = 5'b01111; w[205][76] = 5'b10000; w[205][77] = 5'b00000; w[205][78] = 5'b01111; w[205][79] = 5'b01111; w[205][80] = 5'b00000; w[205][81] = 5'b01111; w[205][82] = 5'b01111; w[205][83] = 5'b01111; w[205][84] = 5'b01111; w[205][85] = 5'b01111; w[205][86] = 5'b01111; w[205][87] = 5'b00000; w[205][88] = 5'b01111; w[205][89] = 5'b01111; w[205][90] = 5'b10000; w[205][91] = 5'b10000; w[205][92] = 5'b01111; w[205][93] = 5'b01111; w[205][94] = 5'b01111; w[205][95] = 5'b01111; w[205][96] = 5'b01111; w[205][97] = 5'b01111; w[205][98] = 5'b01111; w[205][99] = 5'b01111; w[205][100] = 5'b01111; w[205][101] = 5'b00000; w[205][102] = 5'b01111; w[205][103] = 5'b01111; w[205][104] = 5'b10000; w[205][105] = 5'b10000; w[205][106] = 5'b01111; w[205][107] = 5'b00000; w[205][108] = 5'b00000; w[205][109] = 5'b01111; w[205][110] = 5'b01111; w[205][111] = 5'b01111; w[205][112] = 5'b01111; w[205][113] = 5'b01111; w[205][114] = 5'b01111; w[205][115] = 5'b00000; w[205][116] = 5'b01111; w[205][117] = 5'b01111; w[205][118] = 5'b10000; w[205][119] = 5'b10000; w[205][120] = 5'b00000; w[205][121] = 5'b00000; w[205][122] = 5'b00000; w[205][123] = 5'b01111; w[205][124] = 5'b01111; w[205][125] = 5'b01111; w[205][126] = 5'b01111; w[205][127] = 5'b01111; w[205][128] = 5'b01111; w[205][129] = 5'b00000; w[205][130] = 5'b01111; w[205][131] = 5'b01111; w[205][132] = 5'b00000; w[205][133] = 5'b10000; w[205][134] = 5'b01111; w[205][135] = 5'b01111; w[205][136] = 5'b00000; w[205][137] = 5'b01111; w[205][138] = 5'b01111; w[205][139] = 5'b01111; w[205][140] = 5'b01111; w[205][141] = 5'b01111; w[205][142] = 5'b01111; w[205][143] = 5'b00000; w[205][144] = 5'b00000; w[205][145] = 5'b01111; w[205][146] = 5'b00000; w[205][147] = 5'b10000; w[205][148] = 5'b01111; w[205][149] = 5'b00000; w[205][150] = 5'b00000; w[205][151] = 5'b01111; w[205][152] = 5'b01111; w[205][153] = 5'b01111; w[205][154] = 5'b01111; w[205][155] = 5'b01111; w[205][156] = 5'b01111; w[205][157] = 5'b00000; w[205][158] = 5'b00000; w[205][159] = 5'b00000; w[205][160] = 5'b10000; w[205][161] = 5'b10000; w[205][162] = 5'b10000; w[205][163] = 5'b00000; w[205][164] = 5'b00000; w[205][165] = 5'b01111; w[205][166] = 5'b01111; w[205][167] = 5'b01111; w[205][168] = 5'b01111; w[205][169] = 5'b01111; w[205][170] = 5'b01111; w[205][171] = 5'b01111; w[205][172] = 5'b00000; w[205][173] = 5'b00000; w[205][174] = 5'b10000; w[205][175] = 5'b10000; w[205][176] = 5'b10000; w[205][177] = 5'b00000; w[205][178] = 5'b01111; w[205][179] = 5'b01111; w[205][180] = 5'b01111; w[205][181] = 5'b01111; w[205][182] = 5'b01111; w[205][183] = 5'b01111; w[205][184] = 5'b01111; w[205][185] = 5'b01111; w[205][186] = 5'b01111; w[205][187] = 5'b01111; w[205][188] = 5'b01111; w[205][189] = 5'b01111; w[205][190] = 5'b01111; w[205][191] = 5'b01111; w[205][192] = 5'b01111; w[205][193] = 5'b01111; w[205][194] = 5'b01111; w[205][195] = 5'b01111; w[205][196] = 5'b01111; w[205][197] = 5'b01111; w[205][198] = 5'b01111; w[205][199] = 5'b01111; w[205][200] = 5'b01111; w[205][201] = 5'b01111; w[205][202] = 5'b01111; w[205][203] = 5'b01111; w[205][204] = 5'b01111; w[205][205] = 5'b00000; w[205][206] = 5'b01111; w[205][207] = 5'b01111; w[205][208] = 5'b01111; w[205][209] = 5'b01111; 
w[206][0] = 5'b01111; w[206][1] = 5'b01111; w[206][2] = 5'b01111; w[206][3] = 5'b01111; w[206][4] = 5'b01111; w[206][5] = 5'b01111; w[206][6] = 5'b01111; w[206][7] = 5'b01111; w[206][8] = 5'b01111; w[206][9] = 5'b01111; w[206][10] = 5'b01111; w[206][11] = 5'b01111; w[206][12] = 5'b01111; w[206][13] = 5'b01111; w[206][14] = 5'b01111; w[206][15] = 5'b01111; w[206][16] = 5'b01111; w[206][17] = 5'b01111; w[206][18] = 5'b01111; w[206][19] = 5'b01111; w[206][20] = 5'b01111; w[206][21] = 5'b01111; w[206][22] = 5'b01111; w[206][23] = 5'b01111; w[206][24] = 5'b01111; w[206][25] = 5'b01111; w[206][26] = 5'b01111; w[206][27] = 5'b01111; w[206][28] = 5'b01111; w[206][29] = 5'b01111; w[206][30] = 5'b01111; w[206][31] = 5'b00000; w[206][32] = 5'b10000; w[206][33] = 5'b10000; w[206][34] = 5'b10000; w[206][35] = 5'b10000; w[206][36] = 5'b10000; w[206][37] = 5'b10000; w[206][38] = 5'b00000; w[206][39] = 5'b01111; w[206][40] = 5'b01111; w[206][41] = 5'b01111; w[206][42] = 5'b01111; w[206][43] = 5'b01111; w[206][44] = 5'b01111; w[206][45] = 5'b10000; w[206][46] = 5'b10000; w[206][47] = 5'b10000; w[206][48] = 5'b10000; w[206][49] = 5'b10000; w[206][50] = 5'b10000; w[206][51] = 5'b10000; w[206][52] = 5'b10000; w[206][53] = 5'b01111; w[206][54] = 5'b01111; w[206][55] = 5'b01111; w[206][56] = 5'b01111; w[206][57] = 5'b01111; w[206][58] = 5'b01111; w[206][59] = 5'b00000; w[206][60] = 5'b00000; w[206][61] = 5'b01111; w[206][62] = 5'b10000; w[206][63] = 5'b00000; w[206][64] = 5'b01111; w[206][65] = 5'b00000; w[206][66] = 5'b00000; w[206][67] = 5'b01111; w[206][68] = 5'b01111; w[206][69] = 5'b01111; w[206][70] = 5'b01111; w[206][71] = 5'b01111; w[206][72] = 5'b01111; w[206][73] = 5'b00000; w[206][74] = 5'b01111; w[206][75] = 5'b01111; w[206][76] = 5'b10000; w[206][77] = 5'b00000; w[206][78] = 5'b01111; w[206][79] = 5'b01111; w[206][80] = 5'b00000; w[206][81] = 5'b01111; w[206][82] = 5'b01111; w[206][83] = 5'b01111; w[206][84] = 5'b01111; w[206][85] = 5'b01111; w[206][86] = 5'b01111; w[206][87] = 5'b00000; w[206][88] = 5'b01111; w[206][89] = 5'b01111; w[206][90] = 5'b10000; w[206][91] = 5'b10000; w[206][92] = 5'b01111; w[206][93] = 5'b01111; w[206][94] = 5'b01111; w[206][95] = 5'b01111; w[206][96] = 5'b01111; w[206][97] = 5'b01111; w[206][98] = 5'b01111; w[206][99] = 5'b01111; w[206][100] = 5'b01111; w[206][101] = 5'b00000; w[206][102] = 5'b01111; w[206][103] = 5'b01111; w[206][104] = 5'b10000; w[206][105] = 5'b10000; w[206][106] = 5'b01111; w[206][107] = 5'b00000; w[206][108] = 5'b00000; w[206][109] = 5'b01111; w[206][110] = 5'b01111; w[206][111] = 5'b01111; w[206][112] = 5'b01111; w[206][113] = 5'b01111; w[206][114] = 5'b01111; w[206][115] = 5'b00000; w[206][116] = 5'b01111; w[206][117] = 5'b01111; w[206][118] = 5'b10000; w[206][119] = 5'b10000; w[206][120] = 5'b00000; w[206][121] = 5'b00000; w[206][122] = 5'b00000; w[206][123] = 5'b01111; w[206][124] = 5'b01111; w[206][125] = 5'b01111; w[206][126] = 5'b01111; w[206][127] = 5'b01111; w[206][128] = 5'b01111; w[206][129] = 5'b00000; w[206][130] = 5'b01111; w[206][131] = 5'b01111; w[206][132] = 5'b00000; w[206][133] = 5'b10000; w[206][134] = 5'b01111; w[206][135] = 5'b01111; w[206][136] = 5'b00000; w[206][137] = 5'b01111; w[206][138] = 5'b01111; w[206][139] = 5'b01111; w[206][140] = 5'b01111; w[206][141] = 5'b01111; w[206][142] = 5'b01111; w[206][143] = 5'b00000; w[206][144] = 5'b00000; w[206][145] = 5'b01111; w[206][146] = 5'b00000; w[206][147] = 5'b10000; w[206][148] = 5'b01111; w[206][149] = 5'b00000; w[206][150] = 5'b00000; w[206][151] = 5'b01111; w[206][152] = 5'b01111; w[206][153] = 5'b01111; w[206][154] = 5'b01111; w[206][155] = 5'b01111; w[206][156] = 5'b01111; w[206][157] = 5'b00000; w[206][158] = 5'b00000; w[206][159] = 5'b00000; w[206][160] = 5'b10000; w[206][161] = 5'b10000; w[206][162] = 5'b10000; w[206][163] = 5'b00000; w[206][164] = 5'b00000; w[206][165] = 5'b01111; w[206][166] = 5'b01111; w[206][167] = 5'b01111; w[206][168] = 5'b01111; w[206][169] = 5'b01111; w[206][170] = 5'b01111; w[206][171] = 5'b01111; w[206][172] = 5'b00000; w[206][173] = 5'b00000; w[206][174] = 5'b10000; w[206][175] = 5'b10000; w[206][176] = 5'b10000; w[206][177] = 5'b00000; w[206][178] = 5'b01111; w[206][179] = 5'b01111; w[206][180] = 5'b01111; w[206][181] = 5'b01111; w[206][182] = 5'b01111; w[206][183] = 5'b01111; w[206][184] = 5'b01111; w[206][185] = 5'b01111; w[206][186] = 5'b01111; w[206][187] = 5'b01111; w[206][188] = 5'b01111; w[206][189] = 5'b01111; w[206][190] = 5'b01111; w[206][191] = 5'b01111; w[206][192] = 5'b01111; w[206][193] = 5'b01111; w[206][194] = 5'b01111; w[206][195] = 5'b01111; w[206][196] = 5'b01111; w[206][197] = 5'b01111; w[206][198] = 5'b01111; w[206][199] = 5'b01111; w[206][200] = 5'b01111; w[206][201] = 5'b01111; w[206][202] = 5'b01111; w[206][203] = 5'b01111; w[206][204] = 5'b01111; w[206][205] = 5'b01111; w[206][206] = 5'b00000; w[206][207] = 5'b01111; w[206][208] = 5'b01111; w[206][209] = 5'b01111; 
w[207][0] = 5'b01111; w[207][1] = 5'b01111; w[207][2] = 5'b01111; w[207][3] = 5'b01111; w[207][4] = 5'b01111; w[207][5] = 5'b01111; w[207][6] = 5'b01111; w[207][7] = 5'b01111; w[207][8] = 5'b01111; w[207][9] = 5'b01111; w[207][10] = 5'b01111; w[207][11] = 5'b01111; w[207][12] = 5'b01111; w[207][13] = 5'b01111; w[207][14] = 5'b01111; w[207][15] = 5'b01111; w[207][16] = 5'b01111; w[207][17] = 5'b01111; w[207][18] = 5'b01111; w[207][19] = 5'b01111; w[207][20] = 5'b01111; w[207][21] = 5'b01111; w[207][22] = 5'b01111; w[207][23] = 5'b01111; w[207][24] = 5'b01111; w[207][25] = 5'b01111; w[207][26] = 5'b01111; w[207][27] = 5'b01111; w[207][28] = 5'b01111; w[207][29] = 5'b01111; w[207][30] = 5'b01111; w[207][31] = 5'b00000; w[207][32] = 5'b10000; w[207][33] = 5'b10000; w[207][34] = 5'b10000; w[207][35] = 5'b10000; w[207][36] = 5'b10000; w[207][37] = 5'b10000; w[207][38] = 5'b00000; w[207][39] = 5'b01111; w[207][40] = 5'b01111; w[207][41] = 5'b01111; w[207][42] = 5'b01111; w[207][43] = 5'b01111; w[207][44] = 5'b01111; w[207][45] = 5'b10000; w[207][46] = 5'b10000; w[207][47] = 5'b10000; w[207][48] = 5'b10000; w[207][49] = 5'b10000; w[207][50] = 5'b10000; w[207][51] = 5'b10000; w[207][52] = 5'b10000; w[207][53] = 5'b01111; w[207][54] = 5'b01111; w[207][55] = 5'b01111; w[207][56] = 5'b01111; w[207][57] = 5'b01111; w[207][58] = 5'b01111; w[207][59] = 5'b00000; w[207][60] = 5'b00000; w[207][61] = 5'b01111; w[207][62] = 5'b10000; w[207][63] = 5'b00000; w[207][64] = 5'b01111; w[207][65] = 5'b00000; w[207][66] = 5'b00000; w[207][67] = 5'b01111; w[207][68] = 5'b01111; w[207][69] = 5'b01111; w[207][70] = 5'b01111; w[207][71] = 5'b01111; w[207][72] = 5'b01111; w[207][73] = 5'b00000; w[207][74] = 5'b01111; w[207][75] = 5'b01111; w[207][76] = 5'b10000; w[207][77] = 5'b00000; w[207][78] = 5'b01111; w[207][79] = 5'b01111; w[207][80] = 5'b00000; w[207][81] = 5'b01111; w[207][82] = 5'b01111; w[207][83] = 5'b01111; w[207][84] = 5'b01111; w[207][85] = 5'b01111; w[207][86] = 5'b01111; w[207][87] = 5'b00000; w[207][88] = 5'b01111; w[207][89] = 5'b01111; w[207][90] = 5'b10000; w[207][91] = 5'b10000; w[207][92] = 5'b01111; w[207][93] = 5'b01111; w[207][94] = 5'b01111; w[207][95] = 5'b01111; w[207][96] = 5'b01111; w[207][97] = 5'b01111; w[207][98] = 5'b01111; w[207][99] = 5'b01111; w[207][100] = 5'b01111; w[207][101] = 5'b00000; w[207][102] = 5'b01111; w[207][103] = 5'b01111; w[207][104] = 5'b10000; w[207][105] = 5'b10000; w[207][106] = 5'b01111; w[207][107] = 5'b00000; w[207][108] = 5'b00000; w[207][109] = 5'b01111; w[207][110] = 5'b01111; w[207][111] = 5'b01111; w[207][112] = 5'b01111; w[207][113] = 5'b01111; w[207][114] = 5'b01111; w[207][115] = 5'b00000; w[207][116] = 5'b01111; w[207][117] = 5'b01111; w[207][118] = 5'b10000; w[207][119] = 5'b10000; w[207][120] = 5'b00000; w[207][121] = 5'b00000; w[207][122] = 5'b00000; w[207][123] = 5'b01111; w[207][124] = 5'b01111; w[207][125] = 5'b01111; w[207][126] = 5'b01111; w[207][127] = 5'b01111; w[207][128] = 5'b01111; w[207][129] = 5'b00000; w[207][130] = 5'b01111; w[207][131] = 5'b01111; w[207][132] = 5'b00000; w[207][133] = 5'b10000; w[207][134] = 5'b01111; w[207][135] = 5'b01111; w[207][136] = 5'b00000; w[207][137] = 5'b01111; w[207][138] = 5'b01111; w[207][139] = 5'b01111; w[207][140] = 5'b01111; w[207][141] = 5'b01111; w[207][142] = 5'b01111; w[207][143] = 5'b00000; w[207][144] = 5'b00000; w[207][145] = 5'b01111; w[207][146] = 5'b00000; w[207][147] = 5'b10000; w[207][148] = 5'b01111; w[207][149] = 5'b00000; w[207][150] = 5'b00000; w[207][151] = 5'b01111; w[207][152] = 5'b01111; w[207][153] = 5'b01111; w[207][154] = 5'b01111; w[207][155] = 5'b01111; w[207][156] = 5'b01111; w[207][157] = 5'b00000; w[207][158] = 5'b00000; w[207][159] = 5'b00000; w[207][160] = 5'b10000; w[207][161] = 5'b10000; w[207][162] = 5'b10000; w[207][163] = 5'b00000; w[207][164] = 5'b00000; w[207][165] = 5'b01111; w[207][166] = 5'b01111; w[207][167] = 5'b01111; w[207][168] = 5'b01111; w[207][169] = 5'b01111; w[207][170] = 5'b01111; w[207][171] = 5'b01111; w[207][172] = 5'b00000; w[207][173] = 5'b00000; w[207][174] = 5'b10000; w[207][175] = 5'b10000; w[207][176] = 5'b10000; w[207][177] = 5'b00000; w[207][178] = 5'b01111; w[207][179] = 5'b01111; w[207][180] = 5'b01111; w[207][181] = 5'b01111; w[207][182] = 5'b01111; w[207][183] = 5'b01111; w[207][184] = 5'b01111; w[207][185] = 5'b01111; w[207][186] = 5'b01111; w[207][187] = 5'b01111; w[207][188] = 5'b01111; w[207][189] = 5'b01111; w[207][190] = 5'b01111; w[207][191] = 5'b01111; w[207][192] = 5'b01111; w[207][193] = 5'b01111; w[207][194] = 5'b01111; w[207][195] = 5'b01111; w[207][196] = 5'b01111; w[207][197] = 5'b01111; w[207][198] = 5'b01111; w[207][199] = 5'b01111; w[207][200] = 5'b01111; w[207][201] = 5'b01111; w[207][202] = 5'b01111; w[207][203] = 5'b01111; w[207][204] = 5'b01111; w[207][205] = 5'b01111; w[207][206] = 5'b01111; w[207][207] = 5'b00000; w[207][208] = 5'b01111; w[207][209] = 5'b01111; 
w[208][0] = 5'b01111; w[208][1] = 5'b01111; w[208][2] = 5'b01111; w[208][3] = 5'b01111; w[208][4] = 5'b01111; w[208][5] = 5'b01111; w[208][6] = 5'b01111; w[208][7] = 5'b01111; w[208][8] = 5'b01111; w[208][9] = 5'b01111; w[208][10] = 5'b01111; w[208][11] = 5'b01111; w[208][12] = 5'b01111; w[208][13] = 5'b01111; w[208][14] = 5'b01111; w[208][15] = 5'b01111; w[208][16] = 5'b01111; w[208][17] = 5'b01111; w[208][18] = 5'b01111; w[208][19] = 5'b01111; w[208][20] = 5'b01111; w[208][21] = 5'b01111; w[208][22] = 5'b01111; w[208][23] = 5'b01111; w[208][24] = 5'b01111; w[208][25] = 5'b01111; w[208][26] = 5'b01111; w[208][27] = 5'b01111; w[208][28] = 5'b01111; w[208][29] = 5'b01111; w[208][30] = 5'b01111; w[208][31] = 5'b00000; w[208][32] = 5'b10000; w[208][33] = 5'b10000; w[208][34] = 5'b10000; w[208][35] = 5'b10000; w[208][36] = 5'b10000; w[208][37] = 5'b10000; w[208][38] = 5'b00000; w[208][39] = 5'b01111; w[208][40] = 5'b01111; w[208][41] = 5'b01111; w[208][42] = 5'b01111; w[208][43] = 5'b01111; w[208][44] = 5'b01111; w[208][45] = 5'b10000; w[208][46] = 5'b10000; w[208][47] = 5'b10000; w[208][48] = 5'b10000; w[208][49] = 5'b10000; w[208][50] = 5'b10000; w[208][51] = 5'b10000; w[208][52] = 5'b10000; w[208][53] = 5'b01111; w[208][54] = 5'b01111; w[208][55] = 5'b01111; w[208][56] = 5'b01111; w[208][57] = 5'b01111; w[208][58] = 5'b01111; w[208][59] = 5'b00000; w[208][60] = 5'b00000; w[208][61] = 5'b01111; w[208][62] = 5'b10000; w[208][63] = 5'b00000; w[208][64] = 5'b01111; w[208][65] = 5'b00000; w[208][66] = 5'b00000; w[208][67] = 5'b01111; w[208][68] = 5'b01111; w[208][69] = 5'b01111; w[208][70] = 5'b01111; w[208][71] = 5'b01111; w[208][72] = 5'b01111; w[208][73] = 5'b00000; w[208][74] = 5'b01111; w[208][75] = 5'b01111; w[208][76] = 5'b10000; w[208][77] = 5'b00000; w[208][78] = 5'b01111; w[208][79] = 5'b01111; w[208][80] = 5'b00000; w[208][81] = 5'b01111; w[208][82] = 5'b01111; w[208][83] = 5'b01111; w[208][84] = 5'b01111; w[208][85] = 5'b01111; w[208][86] = 5'b01111; w[208][87] = 5'b00000; w[208][88] = 5'b01111; w[208][89] = 5'b01111; w[208][90] = 5'b10000; w[208][91] = 5'b10000; w[208][92] = 5'b01111; w[208][93] = 5'b01111; w[208][94] = 5'b01111; w[208][95] = 5'b01111; w[208][96] = 5'b01111; w[208][97] = 5'b01111; w[208][98] = 5'b01111; w[208][99] = 5'b01111; w[208][100] = 5'b01111; w[208][101] = 5'b00000; w[208][102] = 5'b01111; w[208][103] = 5'b01111; w[208][104] = 5'b10000; w[208][105] = 5'b10000; w[208][106] = 5'b01111; w[208][107] = 5'b00000; w[208][108] = 5'b00000; w[208][109] = 5'b01111; w[208][110] = 5'b01111; w[208][111] = 5'b01111; w[208][112] = 5'b01111; w[208][113] = 5'b01111; w[208][114] = 5'b01111; w[208][115] = 5'b00000; w[208][116] = 5'b01111; w[208][117] = 5'b01111; w[208][118] = 5'b10000; w[208][119] = 5'b10000; w[208][120] = 5'b00000; w[208][121] = 5'b00000; w[208][122] = 5'b00000; w[208][123] = 5'b01111; w[208][124] = 5'b01111; w[208][125] = 5'b01111; w[208][126] = 5'b01111; w[208][127] = 5'b01111; w[208][128] = 5'b01111; w[208][129] = 5'b00000; w[208][130] = 5'b01111; w[208][131] = 5'b01111; w[208][132] = 5'b00000; w[208][133] = 5'b10000; w[208][134] = 5'b01111; w[208][135] = 5'b01111; w[208][136] = 5'b00000; w[208][137] = 5'b01111; w[208][138] = 5'b01111; w[208][139] = 5'b01111; w[208][140] = 5'b01111; w[208][141] = 5'b01111; w[208][142] = 5'b01111; w[208][143] = 5'b00000; w[208][144] = 5'b00000; w[208][145] = 5'b01111; w[208][146] = 5'b00000; w[208][147] = 5'b10000; w[208][148] = 5'b01111; w[208][149] = 5'b00000; w[208][150] = 5'b00000; w[208][151] = 5'b01111; w[208][152] = 5'b01111; w[208][153] = 5'b01111; w[208][154] = 5'b01111; w[208][155] = 5'b01111; w[208][156] = 5'b01111; w[208][157] = 5'b00000; w[208][158] = 5'b00000; w[208][159] = 5'b00000; w[208][160] = 5'b10000; w[208][161] = 5'b10000; w[208][162] = 5'b10000; w[208][163] = 5'b00000; w[208][164] = 5'b00000; w[208][165] = 5'b01111; w[208][166] = 5'b01111; w[208][167] = 5'b01111; w[208][168] = 5'b01111; w[208][169] = 5'b01111; w[208][170] = 5'b01111; w[208][171] = 5'b01111; w[208][172] = 5'b00000; w[208][173] = 5'b00000; w[208][174] = 5'b10000; w[208][175] = 5'b10000; w[208][176] = 5'b10000; w[208][177] = 5'b00000; w[208][178] = 5'b01111; w[208][179] = 5'b01111; w[208][180] = 5'b01111; w[208][181] = 5'b01111; w[208][182] = 5'b01111; w[208][183] = 5'b01111; w[208][184] = 5'b01111; w[208][185] = 5'b01111; w[208][186] = 5'b01111; w[208][187] = 5'b01111; w[208][188] = 5'b01111; w[208][189] = 5'b01111; w[208][190] = 5'b01111; w[208][191] = 5'b01111; w[208][192] = 5'b01111; w[208][193] = 5'b01111; w[208][194] = 5'b01111; w[208][195] = 5'b01111; w[208][196] = 5'b01111; w[208][197] = 5'b01111; w[208][198] = 5'b01111; w[208][199] = 5'b01111; w[208][200] = 5'b01111; w[208][201] = 5'b01111; w[208][202] = 5'b01111; w[208][203] = 5'b01111; w[208][204] = 5'b01111; w[208][205] = 5'b01111; w[208][206] = 5'b01111; w[208][207] = 5'b01111; w[208][208] = 5'b00000; w[208][209] = 5'b01111; 
w[209][0] = 5'b01111; w[209][1] = 5'b01111; w[209][2] = 5'b01111; w[209][3] = 5'b01111; w[209][4] = 5'b01111; w[209][5] = 5'b01111; w[209][6] = 5'b01111; w[209][7] = 5'b01111; w[209][8] = 5'b01111; w[209][9] = 5'b01111; w[209][10] = 5'b01111; w[209][11] = 5'b01111; w[209][12] = 5'b01111; w[209][13] = 5'b01111; w[209][14] = 5'b01111; w[209][15] = 5'b01111; w[209][16] = 5'b01111; w[209][17] = 5'b01111; w[209][18] = 5'b01111; w[209][19] = 5'b01111; w[209][20] = 5'b01111; w[209][21] = 5'b01111; w[209][22] = 5'b01111; w[209][23] = 5'b01111; w[209][24] = 5'b01111; w[209][25] = 5'b01111; w[209][26] = 5'b01111; w[209][27] = 5'b01111; w[209][28] = 5'b01111; w[209][29] = 5'b01111; w[209][30] = 5'b01111; w[209][31] = 5'b00000; w[209][32] = 5'b10000; w[209][33] = 5'b10000; w[209][34] = 5'b10000; w[209][35] = 5'b10000; w[209][36] = 5'b10000; w[209][37] = 5'b10000; w[209][38] = 5'b00000; w[209][39] = 5'b01111; w[209][40] = 5'b01111; w[209][41] = 5'b01111; w[209][42] = 5'b01111; w[209][43] = 5'b01111; w[209][44] = 5'b01111; w[209][45] = 5'b10000; w[209][46] = 5'b10000; w[209][47] = 5'b10000; w[209][48] = 5'b10000; w[209][49] = 5'b10000; w[209][50] = 5'b10000; w[209][51] = 5'b10000; w[209][52] = 5'b10000; w[209][53] = 5'b01111; w[209][54] = 5'b01111; w[209][55] = 5'b01111; w[209][56] = 5'b01111; w[209][57] = 5'b01111; w[209][58] = 5'b01111; w[209][59] = 5'b00000; w[209][60] = 5'b00000; w[209][61] = 5'b01111; w[209][62] = 5'b10000; w[209][63] = 5'b00000; w[209][64] = 5'b01111; w[209][65] = 5'b00000; w[209][66] = 5'b00000; w[209][67] = 5'b01111; w[209][68] = 5'b01111; w[209][69] = 5'b01111; w[209][70] = 5'b01111; w[209][71] = 5'b01111; w[209][72] = 5'b01111; w[209][73] = 5'b00000; w[209][74] = 5'b01111; w[209][75] = 5'b01111; w[209][76] = 5'b10000; w[209][77] = 5'b00000; w[209][78] = 5'b01111; w[209][79] = 5'b01111; w[209][80] = 5'b00000; w[209][81] = 5'b01111; w[209][82] = 5'b01111; w[209][83] = 5'b01111; w[209][84] = 5'b01111; w[209][85] = 5'b01111; w[209][86] = 5'b01111; w[209][87] = 5'b00000; w[209][88] = 5'b01111; w[209][89] = 5'b01111; w[209][90] = 5'b10000; w[209][91] = 5'b10000; w[209][92] = 5'b01111; w[209][93] = 5'b01111; w[209][94] = 5'b01111; w[209][95] = 5'b01111; w[209][96] = 5'b01111; w[209][97] = 5'b01111; w[209][98] = 5'b01111; w[209][99] = 5'b01111; w[209][100] = 5'b01111; w[209][101] = 5'b00000; w[209][102] = 5'b01111; w[209][103] = 5'b01111; w[209][104] = 5'b10000; w[209][105] = 5'b10000; w[209][106] = 5'b01111; w[209][107] = 5'b00000; w[209][108] = 5'b00000; w[209][109] = 5'b01111; w[209][110] = 5'b01111; w[209][111] = 5'b01111; w[209][112] = 5'b01111; w[209][113] = 5'b01111; w[209][114] = 5'b01111; w[209][115] = 5'b00000; w[209][116] = 5'b01111; w[209][117] = 5'b01111; w[209][118] = 5'b10000; w[209][119] = 5'b10000; w[209][120] = 5'b00000; w[209][121] = 5'b00000; w[209][122] = 5'b00000; w[209][123] = 5'b01111; w[209][124] = 5'b01111; w[209][125] = 5'b01111; w[209][126] = 5'b01111; w[209][127] = 5'b01111; w[209][128] = 5'b01111; w[209][129] = 5'b00000; w[209][130] = 5'b01111; w[209][131] = 5'b01111; w[209][132] = 5'b00000; w[209][133] = 5'b10000; w[209][134] = 5'b01111; w[209][135] = 5'b01111; w[209][136] = 5'b00000; w[209][137] = 5'b01111; w[209][138] = 5'b01111; w[209][139] = 5'b01111; w[209][140] = 5'b01111; w[209][141] = 5'b01111; w[209][142] = 5'b01111; w[209][143] = 5'b00000; w[209][144] = 5'b00000; w[209][145] = 5'b01111; w[209][146] = 5'b00000; w[209][147] = 5'b10000; w[209][148] = 5'b01111; w[209][149] = 5'b00000; w[209][150] = 5'b00000; w[209][151] = 5'b01111; w[209][152] = 5'b01111; w[209][153] = 5'b01111; w[209][154] = 5'b01111; w[209][155] = 5'b01111; w[209][156] = 5'b01111; w[209][157] = 5'b00000; w[209][158] = 5'b00000; w[209][159] = 5'b00000; w[209][160] = 5'b10000; w[209][161] = 5'b10000; w[209][162] = 5'b10000; w[209][163] = 5'b00000; w[209][164] = 5'b00000; w[209][165] = 5'b01111; w[209][166] = 5'b01111; w[209][167] = 5'b01111; w[209][168] = 5'b01111; w[209][169] = 5'b01111; w[209][170] = 5'b01111; w[209][171] = 5'b01111; w[209][172] = 5'b00000; w[209][173] = 5'b00000; w[209][174] = 5'b10000; w[209][175] = 5'b10000; w[209][176] = 5'b10000; w[209][177] = 5'b00000; w[209][178] = 5'b01111; w[209][179] = 5'b01111; w[209][180] = 5'b01111; w[209][181] = 5'b01111; w[209][182] = 5'b01111; w[209][183] = 5'b01111; w[209][184] = 5'b01111; w[209][185] = 5'b01111; w[209][186] = 5'b01111; w[209][187] = 5'b01111; w[209][188] = 5'b01111; w[209][189] = 5'b01111; w[209][190] = 5'b01111; w[209][191] = 5'b01111; w[209][192] = 5'b01111; w[209][193] = 5'b01111; w[209][194] = 5'b01111; w[209][195] = 5'b01111; w[209][196] = 5'b01111; w[209][197] = 5'b01111; w[209][198] = 5'b01111; w[209][199] = 5'b01111; w[209][200] = 5'b01111; w[209][201] = 5'b01111; w[209][202] = 5'b01111; w[209][203] = 5'b01111; w[209][204] = 5'b01111; w[209][205] = 5'b01111; w[209][206] = 5'b01111; w[209][207] = 5'b01111; w[209][208] = 5'b01111; w[209][209] = 5'b00000; 
end


    // Generate block for parallel computation of each output n_in[i]
    genvar i, j;
    generate
        for (i = 0; i < n; i = i + 1) begin : synapse_i
            // Array to hold individual terms: w[i][j] * n_out[j]
            wire signed [10:0] term [0:n-1];
            
            // Compute each term based on n_out[j]
            for (j = 0; j < n; j = j + 1) begin : term_j
                assign term[j] = nout[j] ? w[i][j] : -w[i][j];
            end
            
            // Sum all terms combinatorially
//            wire signed [20:0] sum = term[0] + term[1] + term[2] + term[3] + term[4] +
//                                    term[5] + term[6] + term[7] + term[8] + term[9] +
//                                    term[10] + term[11] + term[12] + term[13] + term[14];
               wire signed [20:0] sum = 
                    term[0] + term[1] + term[2] + term[3] + term[4] +
                    term[5] + term[6] + term[7] + term[8] + term[9] +
                    term[10] + term[11] + term[12] + term[13] + term[14] +
                    term[15] + term[16] + term[17] + term[18] + term[19] +
                    term[20] + term[21] + term[22] + term[23] + term[24] +
                    term[25] + term[26] + term[27] + term[28] + term[29] +
                    term[30] + term[31] + term[32] + term[33] + term[34] +
                    term[35] + term[36] + term[37] + term[38] + term[39] +
                    term[40] + term[41] + term[42] + term[43] + term[44] +
                    term[45] + term[46] + term[47] + term[48] + term[49] +
                    term[50] + term[51] + term[52] + term[53] + term[54] +
                    term[55] + term[56] + term[57] + term[58] + term[59] +
                    term[60] + term[61] + term[62] + term[63] + term[64] +
                    term[65] + term[66] + term[67] + term[68] + term[69] +
                    term[70] + term[71] + term[72] + term[73] + term[74] +
                    term[75] + term[76] + term[77] + term[78] + term[79] +
                    term[80] + term[81] + term[82] + term[83] + term[84] +
                    term[85] + term[86] + term[87] + term[88] + term[89] +
                    term[90] + term[91] + term[92] + term[93] + term[94] +
                    term[95] + term[96] + term[97] + term[98] + term[99] +
                    term[100] + term[101] + term[102] + term[103] + term[104] +
                    term[105] + term[106] + term[107] + term[108] + term[109] +
                    term[110] + term[111] + term[112] + term[113] + term[114] +
                    term[115] + term[116] + term[117] + term[118] + term[119] +
                    term[120] + term[121] + term[122] + term[123] + term[124] +
                    term[125] + term[126] + term[127] + term[128] + term[129] +
                    term[130] + term[131] + term[132] + term[133] + term[134] +
                    term[135] + term[136] + term[137] + term[138] + term[139] +
                    term[140] + term[141] + term[142] + term[143] + term[144] +
                    term[145] + term[146] + term[147] + term[148] + term[149] +
                    term[150] + term[151] + term[152] + term[153] + term[154] +
                    term[155] + term[156] + term[157] + term[158] + term[159] +
                    term[160] + term[161] + term[162] + term[163] + term[164] +
                    term[165] + term[166] + term[167] + term[168] + term[169] +
                    term[170] + term[171] + term[172] + term[173] + term[174] +
                    term[175] + term[176] + term[177] + term[178] + term[179] +
                    term[180] + term[181] + term[182] + term[183] + term[184] +
                    term[185] + term[186] + term[187] + term[188] + term[189] +
                    term[190] + term[191] + term[192] + term[193] + term[194] +
                    term[195] + term[196] + term[197] + term[198] + term[199] +
                    term[200] + term[201] + term[202] + term[203] + term[204] +
                    term[205] + term[206] + term[207] + term[208] + term[209] ;
                           

            // Assign n_in[i] based on the sign of the sum
            
            assign nin[i] = (sum > 0) ? 1'b1 : 1'b0;
        end
    endgenerate

endmodule
