`timescale 1ns / 1ps
//module img_load(
//    input [2:0] img_no,
//    input start,
//    input re,
//    input sclk,
//    output reg data_in,
//    output reg load
//);
`timescale 1ns/1ps
module letter_load#(parameter n=210,I=0,T=1,G=2,N=3)(
   input [2:0]img_no,
   input start,
   input re,
   input sclk,
   input [1:0]letter,
   output reg data_in,
   output reg load
    );
reg [0:4*n-1] state;
reg [10:0] c=0;


always @(posedge sclk) begin
        if (re == 1) begin
            load <= 0;
            c <= 0;
            case(letter)
            I:begin
            case(img_no)
            0: state <= 840'h888888888888888888888888888888888100188888888881001888888888880088888888888800888888888888008888888888880088888888888800888888888888008888888888880088888888888100188888888881001888888888888888888888888888888888;
            1: state <= 840'h888888888888888888888888888888888100188888888881331888888888880088888888888800888888888888008888888888880088888888888803888888888888008888888888880088888888888300388888888881301888888888888888888888888888888888;
            2: state <= 840'h884888488848888888884888888888888100188488848881001888448888880088488888888800488888888888008848848888480088488884888800888888888888008488888884880088888888888100188848888881001888884888888888888888884888848888;
            3: state <= 840'h888888888888888888888888888888888180888888888881001888888888880088888888888800888888888888008888888888880888888888888800888888888888808888888888880088888888888100188888888881808888888888888888888888888888888888;
            4: state <= 840'h888808880888888088888888888088888100188888808881001808888888880088888888888800888888888808008888888888880088880880888800888888888888008888888888880080888888088100188808888881001888880888888888088888880888888888;
            5: state <= 840'h888888888288288882888888888888888100588888888881051888828888880588888882888800888888888888008888888888880588888828828800888828888888508882888888880088888888888100188888828881051882888888888888888888888882888888;
            6: state <= 840'h888888808880888888888888888880888808188888888881001888888880888088880888888800888088888888008088888888880088888888888800888888880888008888808088888088808888888100188888888088081888888888888888888088888808888888;
            endcase
            end
            T:begin
            case(img_no)
            0: state <= 840'h888888888888888888888888888888000100100088880001001000888888880088888888888800888888888888008888888888880088888888888800888888888888008888888888880088888888888800888888888888008888888888888888888888888888888888;
            1: state <= 840'h888888888888888888888888888888000300303088880301003000888888880388888888888800888888888888008888888888883088888888888803888888888888008888888888880088888888888803888888888888308888888888888888888888888888888888;
            2: state <= 840'h488884888848888888888888888888000100100088840001001000848888880088888888888800848888488888008888888884880088848888888800848888888884008888488488880088888888888800888888888888008884848884888888888884888848848888;
            3: state <= 840'h888888888888888888888888888888800800800088880001801080888888880088888888888800888888888888008888888888880888888888888800888888888888008888888888880088888888888880888888888888088888888888888888888888888888888888;
            4: state <= 840'h880888088880888088888888880888000100100088880001001000888888880088888888888000888808088888008888888888880088880888888800808888888888008888888880880088888880888800888088888888008888808888888888888880888888088888;
            5: state <= 840'h888288828882888888888888888888050500150088280501001050888888885088888288888800888888882888008288888888880088888888888805888888888288008888282888880088888888888205828888888888508888888828888888828888828888288888;
            6: state <= 840'h808888808888888888888888888888000108100888880808001000888888880088888808888808888808888888008888888088888088888888888800888088888088008888888888888080888088888800888888888888088888888888888888888888088888088888;
            endcase
            end
            G:begin
            case(img_no)
            0: state <= 840'h888888888888888888888888888888880000008888888000000008888800088880008888008888880088880088888888888800888800008888008888000088880088888800888800088880008888800000000888888800000088888888888888888888888888888888;
            1: state <= 840'h888888888888888888888888888888880003008888888030000008888800088880008888038888880388883088888888888800888830008888008888000088883088888830888800388880008888800000000888888803030088888888888888888888888888888888;
            2: state <= 840'h888488884888888888888888888848880000008888888000000008888800088880008484008848880088880048848488888800888800008888008488000084880088888800888800088480008848800000000888888800000088888884888888888488888888888488;
            3: state <= 840'h888888888888888888888888888888880008008888888000000008888808088880808888008888880088880088888888888880888880088888008888000088880088888880888808088880008888800000000888888808000888888888888888888888888888888888;
            4: state <= 840'h088808088888088888888888888880880000008888888000000008808800088080008888008808880088880080808808880800888000008888008880000088880080888800808800088880008888800000000888888800000088888888888888888080888808888888;
            5: state <= 840'h288888288888888888888888828888880505008888888000000008888800088880508888058882280088880028888888882800882850008288508888000088880088288800888800588280058882800000500888888805000088828828888888888888888828828828;
            6: state <= 840'h888808880888880888888888880888080080008888888008000008888880088880808888008888080080880888088888888800888808008888008008008088880888888800800800088880008888800080000888888800008080888088888888888888880888808880;
            endcase
            end
            N:begin
            case(img_no)
            0: state <= 840'h888888888888888888888888888888800088800888888000888008888880000880088888800008800888888000008008888880080080088888800800000888888008800008888880088000088888800888000888888008880008888888888888888888888888888888;
            1: state <= 840'h888888888888888888888888888888803088800888888000888308888880000880088888803008800888888000308008888880080080088888800800003888888008830308888883088000088888800888003888888008883008888888888888888888888888888888;
            2: state <= 840'h848888848884888888888888888888800084800888888000888008848880000880088848800008400888888000008008888880040080088488800800000888888008800008884880048000088888800888000848888008480008888888888888888888488888848888;
            3: state <= 840'h888888888888888888888888888888808088800888888000888088888880000880088888808008800888888000008008888880080880088888808800008888888008808008888880088800088888880888000888888008880808888888888888888888888888888888;
            4: state <= 840'h888888808888800888888880888888800080800888888000888008888080000080088888800008800888888000008008888880080080088888800800000880088000800008888880088000088888800808000888888008800008088088888888888888888888088888;
            5: state <= 840'h888882888888888888888888888888800088800288888050828008888880000880088828800008800888888000558008888885080085088888800800000888888008800008828880088000588888805288500888888008880008888288888888888888888888288888;
            6: state <= 840'h888888088888888888888888888808800088808808888000808008888880800880088888800008800888888000008088888880080080088888880808000888888008800008888880088000888888808088000888808008880808888888880888888888888888888808;            
            endcase
            end    
        endcase
        end
        else if (start == 1) begin
            if (c <(4*n)) begin
                load <= 1;
                data_in <= state[4*n-1];         // Send MSB first
                state <= state >> 1;          // Left shift by 1
                c <= c + 1;
            end
            else begin
                load <= 0;
            end
        end
        else begin
            load <= 0;
        end
    end

endmodule
